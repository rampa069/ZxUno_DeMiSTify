
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e4",x"ec",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e4",x"ec",x"c2"),
    14 => (x"48",x"f4",x"d9",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e4",x"dc"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"48",x"72",x"4c"),
    72 => (x"7c",x"70",x"98",x"ff"),
    73 => (x"bf",x"f4",x"d9",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"ff",x"c3",x"48",x"71"),
    79 => (x"d0",x"7c",x"70",x"98"),
    80 => (x"29",x"d0",x"49",x"66"),
    81 => (x"ff",x"c3",x"48",x"71"),
    82 => (x"d0",x"7c",x"70",x"98"),
    83 => (x"29",x"c8",x"49",x"66"),
    84 => (x"ff",x"c3",x"48",x"71"),
    85 => (x"d0",x"7c",x"70",x"98"),
    86 => (x"ff",x"c3",x"48",x"66"),
    87 => (x"72",x"7c",x"70",x"98"),
    88 => (x"71",x"29",x"d0",x"49"),
    89 => (x"98",x"ff",x"c3",x"48"),
    90 => (x"4b",x"6c",x"7c",x"70"),
    91 => (x"4d",x"ff",x"f0",x"c9"),
    92 => (x"05",x"ab",x"ff",x"c3"),
    93 => (x"ff",x"c3",x"87",x"d0"),
    94 => (x"c1",x"4b",x"6c",x"7c"),
    95 => (x"87",x"c6",x"02",x"8d"),
    96 => (x"02",x"ab",x"ff",x"c3"),
    97 => (x"48",x"73",x"87",x"f0"),
    98 => (x"1e",x"87",x"ff",x"fd"),
    99 => (x"d4",x"ff",x"49",x"c0"),
   100 => (x"78",x"ff",x"c3",x"48"),
   101 => (x"c8",x"c3",x"81",x"c1"),
   102 => (x"f1",x"04",x"a9",x"b7"),
   103 => (x"1e",x"4f",x"26",x"87"),
   104 => (x"87",x"e7",x"1e",x"73"),
   105 => (x"4b",x"df",x"f8",x"c4"),
   106 => (x"ff",x"c0",x"1e",x"c0"),
   107 => (x"49",x"f7",x"c1",x"f0"),
   108 => (x"c4",x"87",x"df",x"fd"),
   109 => (x"05",x"a8",x"c1",x"86"),
   110 => (x"ff",x"87",x"ea",x"c0"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c0",x"c0",x"c1",x"78"),
   113 => (x"1e",x"c0",x"c0",x"c0"),
   114 => (x"c1",x"f0",x"e1",x"c0"),
   115 => (x"c1",x"fd",x"49",x"e9"),
   116 => (x"70",x"86",x"c4",x"87"),
   117 => (x"87",x"ca",x"05",x"98"),
   118 => (x"c3",x"48",x"d4",x"ff"),
   119 => (x"48",x"c1",x"78",x"ff"),
   120 => (x"e6",x"fe",x"87",x"cb"),
   121 => (x"05",x"8b",x"c1",x"87"),
   122 => (x"c0",x"87",x"fd",x"fe"),
   123 => (x"87",x"de",x"fc",x"48"),
   124 => (x"ff",x"1e",x"73",x"1e"),
   125 => (x"ff",x"c3",x"48",x"d4"),
   126 => (x"c0",x"4b",x"d3",x"78"),
   127 => (x"f0",x"ff",x"c0",x"1e"),
   128 => (x"fc",x"49",x"c1",x"c1"),
   129 => (x"86",x"c4",x"87",x"cc"),
   130 => (x"ca",x"05",x"98",x"70"),
   131 => (x"48",x"d4",x"ff",x"87"),
   132 => (x"c1",x"78",x"ff",x"c3"),
   133 => (x"fd",x"87",x"cb",x"48"),
   134 => (x"8b",x"c1",x"87",x"f1"),
   135 => (x"87",x"db",x"ff",x"05"),
   136 => (x"e9",x"fb",x"48",x"c0"),
   137 => (x"5b",x"5e",x"0e",x"87"),
   138 => (x"d4",x"ff",x"0e",x"5c"),
   139 => (x"87",x"db",x"fd",x"4c"),
   140 => (x"c0",x"1e",x"ea",x"c6"),
   141 => (x"c8",x"c1",x"f0",x"e1"),
   142 => (x"87",x"d6",x"fb",x"49"),
   143 => (x"a8",x"c1",x"86",x"c4"),
   144 => (x"fe",x"87",x"c8",x"02"),
   145 => (x"48",x"c0",x"87",x"ea"),
   146 => (x"fa",x"87",x"e2",x"c1"),
   147 => (x"49",x"70",x"87",x"d2"),
   148 => (x"99",x"ff",x"ff",x"cf"),
   149 => (x"02",x"a9",x"ea",x"c6"),
   150 => (x"d3",x"fe",x"87",x"c8"),
   151 => (x"c1",x"48",x"c0",x"87"),
   152 => (x"ff",x"c3",x"87",x"cb"),
   153 => (x"4b",x"f1",x"c0",x"7c"),
   154 => (x"70",x"87",x"f4",x"fc"),
   155 => (x"eb",x"c0",x"02",x"98"),
   156 => (x"c0",x"1e",x"c0",x"87"),
   157 => (x"fa",x"c1",x"f0",x"ff"),
   158 => (x"87",x"d6",x"fa",x"49"),
   159 => (x"98",x"70",x"86",x"c4"),
   160 => (x"c3",x"87",x"d9",x"05"),
   161 => (x"49",x"6c",x"7c",x"ff"),
   162 => (x"7c",x"7c",x"ff",x"c3"),
   163 => (x"c0",x"c1",x"7c",x"7c"),
   164 => (x"87",x"c4",x"02",x"99"),
   165 => (x"87",x"d5",x"48",x"c1"),
   166 => (x"87",x"d1",x"48",x"c0"),
   167 => (x"c4",x"05",x"ab",x"c2"),
   168 => (x"c8",x"48",x"c0",x"87"),
   169 => (x"05",x"8b",x"c1",x"87"),
   170 => (x"c0",x"87",x"fd",x"fe"),
   171 => (x"87",x"dc",x"f9",x"48"),
   172 => (x"c2",x"1e",x"73",x"1e"),
   173 => (x"c1",x"48",x"f4",x"d9"),
   174 => (x"ff",x"4b",x"c7",x"78"),
   175 => (x"78",x"c2",x"48",x"d0"),
   176 => (x"ff",x"87",x"c8",x"fb"),
   177 => (x"78",x"c3",x"48",x"d0"),
   178 => (x"e5",x"c0",x"1e",x"c0"),
   179 => (x"49",x"c0",x"c1",x"d0"),
   180 => (x"c4",x"87",x"ff",x"f8"),
   181 => (x"05",x"a8",x"c1",x"86"),
   182 => (x"c2",x"4b",x"87",x"c1"),
   183 => (x"87",x"c5",x"05",x"ab"),
   184 => (x"f9",x"c0",x"48",x"c0"),
   185 => (x"05",x"8b",x"c1",x"87"),
   186 => (x"fc",x"87",x"d0",x"ff"),
   187 => (x"d9",x"c2",x"87",x"f7"),
   188 => (x"98",x"70",x"58",x"f8"),
   189 => (x"c1",x"87",x"cd",x"05"),
   190 => (x"f0",x"ff",x"c0",x"1e"),
   191 => (x"f8",x"49",x"d0",x"c1"),
   192 => (x"86",x"c4",x"87",x"d0"),
   193 => (x"c3",x"48",x"d4",x"ff"),
   194 => (x"fd",x"c2",x"78",x"ff"),
   195 => (x"fc",x"d9",x"c2",x"87"),
   196 => (x"48",x"d0",x"ff",x"58"),
   197 => (x"d4",x"ff",x"78",x"c2"),
   198 => (x"78",x"ff",x"c3",x"48"),
   199 => (x"ed",x"f7",x"48",x"c1"),
   200 => (x"5b",x"5e",x"0e",x"87"),
   201 => (x"71",x"0e",x"5d",x"5c"),
   202 => (x"c5",x"4c",x"c0",x"4b"),
   203 => (x"4a",x"df",x"cd",x"ee"),
   204 => (x"c3",x"48",x"d4",x"ff"),
   205 => (x"48",x"68",x"78",x"ff"),
   206 => (x"05",x"a8",x"fe",x"c3"),
   207 => (x"ff",x"87",x"fe",x"c0"),
   208 => (x"9b",x"73",x"4d",x"d4"),
   209 => (x"d0",x"87",x"cc",x"02"),
   210 => (x"49",x"73",x"1e",x"66"),
   211 => (x"c4",x"87",x"e8",x"f5"),
   212 => (x"ff",x"87",x"d6",x"86"),
   213 => (x"d1",x"c4",x"48",x"d0"),
   214 => (x"7d",x"ff",x"c3",x"78"),
   215 => (x"c1",x"48",x"66",x"d0"),
   216 => (x"58",x"a6",x"d4",x"88"),
   217 => (x"f0",x"05",x"98",x"70"),
   218 => (x"48",x"d4",x"ff",x"87"),
   219 => (x"78",x"78",x"ff",x"c3"),
   220 => (x"c5",x"05",x"9b",x"73"),
   221 => (x"48",x"d0",x"ff",x"87"),
   222 => (x"4a",x"c1",x"78",x"d0"),
   223 => (x"05",x"8a",x"c1",x"4c"),
   224 => (x"74",x"87",x"ed",x"fe"),
   225 => (x"87",x"c2",x"f6",x"48"),
   226 => (x"71",x"1e",x"73",x"1e"),
   227 => (x"ff",x"4b",x"c0",x"4a"),
   228 => (x"ff",x"c3",x"48",x"d4"),
   229 => (x"48",x"d0",x"ff",x"78"),
   230 => (x"ff",x"78",x"c3",x"c4"),
   231 => (x"ff",x"c3",x"48",x"d4"),
   232 => (x"c0",x"1e",x"72",x"78"),
   233 => (x"d1",x"c1",x"f0",x"ff"),
   234 => (x"87",x"e6",x"f5",x"49"),
   235 => (x"98",x"70",x"86",x"c4"),
   236 => (x"c8",x"87",x"d2",x"05"),
   237 => (x"66",x"cc",x"1e",x"c0"),
   238 => (x"87",x"e5",x"fd",x"49"),
   239 => (x"4b",x"70",x"86",x"c4"),
   240 => (x"c2",x"48",x"d0",x"ff"),
   241 => (x"f5",x"48",x"73",x"78"),
   242 => (x"5e",x"0e",x"87",x"c4"),
   243 => (x"0e",x"5d",x"5c",x"5b"),
   244 => (x"ff",x"c0",x"1e",x"c0"),
   245 => (x"49",x"c9",x"c1",x"f0"),
   246 => (x"d2",x"87",x"f7",x"f4"),
   247 => (x"fc",x"d9",x"c2",x"1e"),
   248 => (x"87",x"fd",x"fc",x"49"),
   249 => (x"4c",x"c0",x"86",x"c8"),
   250 => (x"b7",x"d2",x"84",x"c1"),
   251 => (x"87",x"f8",x"04",x"ac"),
   252 => (x"97",x"fc",x"d9",x"c2"),
   253 => (x"c0",x"c3",x"49",x"bf"),
   254 => (x"a9",x"c0",x"c1",x"99"),
   255 => (x"87",x"e7",x"c0",x"05"),
   256 => (x"97",x"c3",x"da",x"c2"),
   257 => (x"31",x"d0",x"49",x"bf"),
   258 => (x"97",x"c4",x"da",x"c2"),
   259 => (x"32",x"c8",x"4a",x"bf"),
   260 => (x"da",x"c2",x"b1",x"72"),
   261 => (x"4a",x"bf",x"97",x"c5"),
   262 => (x"cf",x"4c",x"71",x"b1"),
   263 => (x"9c",x"ff",x"ff",x"ff"),
   264 => (x"34",x"ca",x"84",x"c1"),
   265 => (x"c2",x"87",x"e7",x"c1"),
   266 => (x"bf",x"97",x"c5",x"da"),
   267 => (x"c6",x"31",x"c1",x"49"),
   268 => (x"c6",x"da",x"c2",x"99"),
   269 => (x"c7",x"4a",x"bf",x"97"),
   270 => (x"b1",x"72",x"2a",x"b7"),
   271 => (x"97",x"c1",x"da",x"c2"),
   272 => (x"cf",x"4d",x"4a",x"bf"),
   273 => (x"c2",x"da",x"c2",x"9d"),
   274 => (x"c3",x"4a",x"bf",x"97"),
   275 => (x"c2",x"32",x"ca",x"9a"),
   276 => (x"bf",x"97",x"c3",x"da"),
   277 => (x"73",x"33",x"c2",x"4b"),
   278 => (x"c4",x"da",x"c2",x"b2"),
   279 => (x"c3",x"4b",x"bf",x"97"),
   280 => (x"b7",x"c6",x"9b",x"c0"),
   281 => (x"c2",x"b2",x"73",x"2b"),
   282 => (x"71",x"48",x"c1",x"81"),
   283 => (x"c1",x"49",x"70",x"30"),
   284 => (x"70",x"30",x"75",x"48"),
   285 => (x"c1",x"4c",x"72",x"4d"),
   286 => (x"c8",x"94",x"71",x"84"),
   287 => (x"06",x"ad",x"b7",x"c0"),
   288 => (x"34",x"c1",x"87",x"cc"),
   289 => (x"c0",x"c8",x"2d",x"b7"),
   290 => (x"ff",x"01",x"ad",x"b7"),
   291 => (x"48",x"74",x"87",x"f4"),
   292 => (x"0e",x"87",x"f7",x"f1"),
   293 => (x"5d",x"5c",x"5b",x"5e"),
   294 => (x"c2",x"86",x"f8",x"0e"),
   295 => (x"c0",x"48",x"e2",x"e2"),
   296 => (x"da",x"da",x"c2",x"78"),
   297 => (x"fb",x"49",x"c0",x"1e"),
   298 => (x"86",x"c4",x"87",x"de"),
   299 => (x"c5",x"05",x"98",x"70"),
   300 => (x"c9",x"48",x"c0",x"87"),
   301 => (x"4d",x"c0",x"87",x"c0"),
   302 => (x"ed",x"c0",x"7e",x"c1"),
   303 => (x"c2",x"49",x"bf",x"e6"),
   304 => (x"71",x"4a",x"d0",x"db"),
   305 => (x"e0",x"ee",x"4b",x"c8"),
   306 => (x"05",x"98",x"70",x"87"),
   307 => (x"7e",x"c0",x"87",x"c2"),
   308 => (x"bf",x"e2",x"ed",x"c0"),
   309 => (x"ec",x"db",x"c2",x"49"),
   310 => (x"4b",x"c8",x"71",x"4a"),
   311 => (x"70",x"87",x"ca",x"ee"),
   312 => (x"87",x"c2",x"05",x"98"),
   313 => (x"02",x"6e",x"7e",x"c0"),
   314 => (x"c2",x"87",x"fd",x"c0"),
   315 => (x"4d",x"bf",x"e0",x"e1"),
   316 => (x"9f",x"d8",x"e2",x"c2"),
   317 => (x"c5",x"48",x"7e",x"bf"),
   318 => (x"05",x"a8",x"ea",x"d6"),
   319 => (x"e1",x"c2",x"87",x"c7"),
   320 => (x"ce",x"4d",x"bf",x"e0"),
   321 => (x"ca",x"48",x"6e",x"87"),
   322 => (x"02",x"a8",x"d5",x"e9"),
   323 => (x"48",x"c0",x"87",x"c5"),
   324 => (x"c2",x"87",x"e3",x"c7"),
   325 => (x"75",x"1e",x"da",x"da"),
   326 => (x"87",x"ec",x"f9",x"49"),
   327 => (x"98",x"70",x"86",x"c4"),
   328 => (x"c0",x"87",x"c5",x"05"),
   329 => (x"87",x"ce",x"c7",x"48"),
   330 => (x"bf",x"e2",x"ed",x"c0"),
   331 => (x"ec",x"db",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f2",x"ec"),
   334 => (x"87",x"c8",x"05",x"98"),
   335 => (x"48",x"e2",x"e2",x"c2"),
   336 => (x"87",x"da",x"78",x"c1"),
   337 => (x"bf",x"e6",x"ed",x"c0"),
   338 => (x"d0",x"db",x"c2",x"49"),
   339 => (x"4b",x"c8",x"71",x"4a"),
   340 => (x"70",x"87",x"d6",x"ec"),
   341 => (x"c5",x"c0",x"02",x"98"),
   342 => (x"c6",x"48",x"c0",x"87"),
   343 => (x"e2",x"c2",x"87",x"d8"),
   344 => (x"49",x"bf",x"97",x"d8"),
   345 => (x"05",x"a9",x"d5",x"c1"),
   346 => (x"c2",x"87",x"cd",x"c0"),
   347 => (x"bf",x"97",x"d9",x"e2"),
   348 => (x"a9",x"ea",x"c2",x"49"),
   349 => (x"87",x"c5",x"c0",x"02"),
   350 => (x"f9",x"c5",x"48",x"c0"),
   351 => (x"da",x"da",x"c2",x"87"),
   352 => (x"48",x"7e",x"bf",x"97"),
   353 => (x"02",x"a8",x"e9",x"c3"),
   354 => (x"6e",x"87",x"ce",x"c0"),
   355 => (x"a8",x"eb",x"c3",x"48"),
   356 => (x"87",x"c5",x"c0",x"02"),
   357 => (x"dd",x"c5",x"48",x"c0"),
   358 => (x"e5",x"da",x"c2",x"87"),
   359 => (x"99",x"49",x"bf",x"97"),
   360 => (x"87",x"cc",x"c0",x"05"),
   361 => (x"97",x"e6",x"da",x"c2"),
   362 => (x"a9",x"c2",x"49",x"bf"),
   363 => (x"87",x"c5",x"c0",x"02"),
   364 => (x"c1",x"c5",x"48",x"c0"),
   365 => (x"e7",x"da",x"c2",x"87"),
   366 => (x"c2",x"48",x"bf",x"97"),
   367 => (x"70",x"58",x"de",x"e2"),
   368 => (x"88",x"c1",x"48",x"4c"),
   369 => (x"58",x"e2",x"e2",x"c2"),
   370 => (x"97",x"e8",x"da",x"c2"),
   371 => (x"81",x"75",x"49",x"bf"),
   372 => (x"97",x"e9",x"da",x"c2"),
   373 => (x"32",x"c8",x"4a",x"bf"),
   374 => (x"c2",x"7e",x"a1",x"72"),
   375 => (x"6e",x"48",x"ef",x"e6"),
   376 => (x"ea",x"da",x"c2",x"78"),
   377 => (x"c8",x"48",x"bf",x"97"),
   378 => (x"e2",x"c2",x"58",x"a6"),
   379 => (x"c2",x"02",x"bf",x"e2"),
   380 => (x"ed",x"c0",x"87",x"cf"),
   381 => (x"c2",x"49",x"bf",x"e2"),
   382 => (x"71",x"4a",x"ec",x"db"),
   383 => (x"e8",x"e9",x"4b",x"c8"),
   384 => (x"02",x"98",x"70",x"87"),
   385 => (x"c0",x"87",x"c5",x"c0"),
   386 => (x"87",x"ea",x"c3",x"48"),
   387 => (x"bf",x"da",x"e2",x"c2"),
   388 => (x"c3",x"e7",x"c2",x"4c"),
   389 => (x"ff",x"da",x"c2",x"5c"),
   390 => (x"c8",x"49",x"bf",x"97"),
   391 => (x"fe",x"da",x"c2",x"31"),
   392 => (x"a1",x"4a",x"bf",x"97"),
   393 => (x"c0",x"db",x"c2",x"49"),
   394 => (x"d0",x"4a",x"bf",x"97"),
   395 => (x"49",x"a1",x"72",x"32"),
   396 => (x"97",x"c1",x"db",x"c2"),
   397 => (x"32",x"d8",x"4a",x"bf"),
   398 => (x"c4",x"49",x"a1",x"72"),
   399 => (x"e6",x"c2",x"91",x"66"),
   400 => (x"c2",x"81",x"bf",x"ef"),
   401 => (x"c2",x"59",x"f7",x"e6"),
   402 => (x"bf",x"97",x"c7",x"db"),
   403 => (x"c2",x"32",x"c8",x"4a"),
   404 => (x"bf",x"97",x"c6",x"db"),
   405 => (x"c2",x"4a",x"a2",x"4b"),
   406 => (x"bf",x"97",x"c8",x"db"),
   407 => (x"73",x"33",x"d0",x"4b"),
   408 => (x"db",x"c2",x"4a",x"a2"),
   409 => (x"4b",x"bf",x"97",x"c9"),
   410 => (x"33",x"d8",x"9b",x"cf"),
   411 => (x"c2",x"4a",x"a2",x"73"),
   412 => (x"c2",x"5a",x"fb",x"e6"),
   413 => (x"c2",x"92",x"74",x"8a"),
   414 => (x"72",x"48",x"fb",x"e6"),
   415 => (x"c1",x"c1",x"78",x"a1"),
   416 => (x"ec",x"da",x"c2",x"87"),
   417 => (x"c8",x"49",x"bf",x"97"),
   418 => (x"eb",x"da",x"c2",x"31"),
   419 => (x"a1",x"4a",x"bf",x"97"),
   420 => (x"c7",x"31",x"c5",x"49"),
   421 => (x"29",x"c9",x"81",x"ff"),
   422 => (x"59",x"c3",x"e7",x"c2"),
   423 => (x"97",x"f1",x"da",x"c2"),
   424 => (x"32",x"c8",x"4a",x"bf"),
   425 => (x"97",x"f0",x"da",x"c2"),
   426 => (x"4a",x"a2",x"4b",x"bf"),
   427 => (x"6e",x"92",x"66",x"c4"),
   428 => (x"ff",x"e6",x"c2",x"82"),
   429 => (x"f7",x"e6",x"c2",x"5a"),
   430 => (x"c2",x"78",x"c0",x"48"),
   431 => (x"72",x"48",x"f3",x"e6"),
   432 => (x"e7",x"c2",x"78",x"a1"),
   433 => (x"e6",x"c2",x"48",x"c3"),
   434 => (x"c2",x"78",x"bf",x"f7"),
   435 => (x"c2",x"48",x"c7",x"e7"),
   436 => (x"78",x"bf",x"fb",x"e6"),
   437 => (x"bf",x"e2",x"e2",x"c2"),
   438 => (x"87",x"c9",x"c0",x"02"),
   439 => (x"30",x"c4",x"48",x"74"),
   440 => (x"c9",x"c0",x"7e",x"70"),
   441 => (x"ff",x"e6",x"c2",x"87"),
   442 => (x"30",x"c4",x"48",x"bf"),
   443 => (x"e2",x"c2",x"7e",x"70"),
   444 => (x"78",x"6e",x"48",x"e6"),
   445 => (x"8e",x"f8",x"48",x"c1"),
   446 => (x"4c",x"26",x"4d",x"26"),
   447 => (x"4f",x"26",x"4b",x"26"),
   448 => (x"5c",x"5b",x"5e",x"0e"),
   449 => (x"4a",x"71",x"0e",x"5d"),
   450 => (x"bf",x"e2",x"e2",x"c2"),
   451 => (x"72",x"87",x"cb",x"02"),
   452 => (x"72",x"2b",x"c7",x"4b"),
   453 => (x"9d",x"ff",x"c1",x"4d"),
   454 => (x"4b",x"72",x"87",x"c9"),
   455 => (x"4d",x"72",x"2b",x"c8"),
   456 => (x"c2",x"9d",x"ff",x"c3"),
   457 => (x"83",x"bf",x"ef",x"e6"),
   458 => (x"bf",x"de",x"ed",x"c0"),
   459 => (x"87",x"d9",x"02",x"ab"),
   460 => (x"5b",x"e2",x"ed",x"c0"),
   461 => (x"1e",x"da",x"da",x"c2"),
   462 => (x"cb",x"f1",x"49",x"73"),
   463 => (x"70",x"86",x"c4",x"87"),
   464 => (x"87",x"c5",x"05",x"98"),
   465 => (x"e6",x"c0",x"48",x"c0"),
   466 => (x"e2",x"e2",x"c2",x"87"),
   467 => (x"87",x"d2",x"02",x"bf"),
   468 => (x"91",x"c4",x"49",x"75"),
   469 => (x"81",x"da",x"da",x"c2"),
   470 => (x"ff",x"cf",x"4c",x"69"),
   471 => (x"9c",x"ff",x"ff",x"ff"),
   472 => (x"49",x"75",x"87",x"cb"),
   473 => (x"da",x"c2",x"91",x"c2"),
   474 => (x"69",x"9f",x"81",x"da"),
   475 => (x"fe",x"48",x"74",x"4c"),
   476 => (x"5e",x"0e",x"87",x"c6"),
   477 => (x"0e",x"5d",x"5c",x"5b"),
   478 => (x"4c",x"71",x"86",x"f8"),
   479 => (x"87",x"c5",x"05",x"9c"),
   480 => (x"c0",x"c3",x"48",x"c0"),
   481 => (x"7e",x"a4",x"c8",x"87"),
   482 => (x"d8",x"78",x"c0",x"48"),
   483 => (x"87",x"c7",x"02",x"66"),
   484 => (x"bf",x"97",x"66",x"d8"),
   485 => (x"c0",x"87",x"c5",x"05"),
   486 => (x"87",x"e9",x"c2",x"48"),
   487 => (x"49",x"c1",x"1e",x"c0"),
   488 => (x"87",x"e3",x"c7",x"49"),
   489 => (x"4d",x"70",x"86",x"c4"),
   490 => (x"c2",x"c1",x"02",x"9d"),
   491 => (x"ea",x"e2",x"c2",x"87"),
   492 => (x"49",x"66",x"d8",x"4a"),
   493 => (x"70",x"87",x"d7",x"e2"),
   494 => (x"f2",x"c0",x"02",x"98"),
   495 => (x"d8",x"4a",x"75",x"87"),
   496 => (x"4b",x"cb",x"49",x"66"),
   497 => (x"70",x"87",x"fc",x"e2"),
   498 => (x"e2",x"c0",x"02",x"98"),
   499 => (x"75",x"1e",x"c0",x"87"),
   500 => (x"87",x"c7",x"02",x"9d"),
   501 => (x"c0",x"48",x"a6",x"c8"),
   502 => (x"c8",x"87",x"c5",x"78"),
   503 => (x"78",x"c1",x"48",x"a6"),
   504 => (x"c6",x"49",x"66",x"c8"),
   505 => (x"86",x"c4",x"87",x"e1"),
   506 => (x"05",x"9d",x"4d",x"70"),
   507 => (x"75",x"87",x"fe",x"fe"),
   508 => (x"ce",x"c1",x"02",x"9d"),
   509 => (x"49",x"a5",x"dc",x"87"),
   510 => (x"78",x"69",x"48",x"6e"),
   511 => (x"c4",x"49",x"a5",x"da"),
   512 => (x"a4",x"c4",x"48",x"a6"),
   513 => (x"48",x"69",x"9f",x"78"),
   514 => (x"78",x"08",x"66",x"c4"),
   515 => (x"bf",x"e2",x"e2",x"c2"),
   516 => (x"d4",x"87",x"d2",x"02"),
   517 => (x"69",x"9f",x"49",x"a5"),
   518 => (x"ff",x"ff",x"c0",x"49"),
   519 => (x"d0",x"48",x"71",x"99"),
   520 => (x"c2",x"7e",x"70",x"30"),
   521 => (x"6e",x"7e",x"c0",x"87"),
   522 => (x"bf",x"66",x"c4",x"48"),
   523 => (x"08",x"66",x"c4",x"80"),
   524 => (x"cc",x"7c",x"c0",x"78"),
   525 => (x"66",x"c4",x"49",x"a4"),
   526 => (x"a4",x"d0",x"79",x"bf"),
   527 => (x"c1",x"79",x"c0",x"49"),
   528 => (x"c0",x"87",x"c2",x"48"),
   529 => (x"fa",x"8e",x"f8",x"48"),
   530 => (x"5e",x"0e",x"87",x"ee"),
   531 => (x"71",x"0e",x"5c",x"5b"),
   532 => (x"c1",x"02",x"9c",x"4c"),
   533 => (x"a4",x"c8",x"87",x"cb"),
   534 => (x"c1",x"02",x"69",x"49"),
   535 => (x"49",x"6c",x"87",x"c3"),
   536 => (x"71",x"48",x"66",x"cc"),
   537 => (x"58",x"a6",x"d0",x"80"),
   538 => (x"e2",x"c2",x"b9",x"70"),
   539 => (x"ff",x"4a",x"bf",x"de"),
   540 => (x"71",x"99",x"72",x"ba"),
   541 => (x"e5",x"c0",x"02",x"99"),
   542 => (x"4b",x"a4",x"c4",x"87"),
   543 => (x"ff",x"f9",x"49",x"6b"),
   544 => (x"c2",x"7b",x"70",x"87"),
   545 => (x"49",x"bf",x"da",x"e2"),
   546 => (x"7c",x"71",x"81",x"6c"),
   547 => (x"c2",x"b9",x"66",x"cc"),
   548 => (x"4a",x"bf",x"de",x"e2"),
   549 => (x"99",x"72",x"ba",x"ff"),
   550 => (x"ff",x"05",x"99",x"71"),
   551 => (x"66",x"cc",x"87",x"db"),
   552 => (x"87",x"d6",x"f9",x"7c"),
   553 => (x"71",x"1e",x"73",x"1e"),
   554 => (x"c7",x"02",x"9b",x"4b"),
   555 => (x"49",x"a3",x"c8",x"87"),
   556 => (x"87",x"c5",x"05",x"69"),
   557 => (x"f6",x"c0",x"48",x"c0"),
   558 => (x"f3",x"e6",x"c2",x"87"),
   559 => (x"a3",x"c4",x"49",x"bf"),
   560 => (x"c2",x"4a",x"6a",x"4a"),
   561 => (x"da",x"e2",x"c2",x"8a"),
   562 => (x"a1",x"72",x"92",x"bf"),
   563 => (x"de",x"e2",x"c2",x"49"),
   564 => (x"9a",x"6b",x"4a",x"bf"),
   565 => (x"c0",x"49",x"a1",x"72"),
   566 => (x"c8",x"59",x"e2",x"ed"),
   567 => (x"ea",x"71",x"1e",x"66"),
   568 => (x"86",x"c4",x"87",x"e6"),
   569 => (x"c4",x"05",x"98",x"70"),
   570 => (x"c2",x"48",x"c0",x"87"),
   571 => (x"f8",x"48",x"c1",x"87"),
   572 => (x"73",x"1e",x"87",x"ca"),
   573 => (x"9b",x"4b",x"71",x"1e"),
   574 => (x"87",x"e4",x"c0",x"02"),
   575 => (x"5b",x"c7",x"e7",x"c2"),
   576 => (x"8a",x"c2",x"4a",x"73"),
   577 => (x"bf",x"da",x"e2",x"c2"),
   578 => (x"e6",x"c2",x"92",x"49"),
   579 => (x"72",x"48",x"bf",x"f3"),
   580 => (x"cb",x"e7",x"c2",x"80"),
   581 => (x"c4",x"48",x"71",x"58"),
   582 => (x"ea",x"e2",x"c2",x"30"),
   583 => (x"87",x"ed",x"c0",x"58"),
   584 => (x"48",x"c3",x"e7",x"c2"),
   585 => (x"bf",x"f7",x"e6",x"c2"),
   586 => (x"c7",x"e7",x"c2",x"78"),
   587 => (x"fb",x"e6",x"c2",x"48"),
   588 => (x"e2",x"c2",x"78",x"bf"),
   589 => (x"c9",x"02",x"bf",x"e2"),
   590 => (x"da",x"e2",x"c2",x"87"),
   591 => (x"31",x"c4",x"49",x"bf"),
   592 => (x"e6",x"c2",x"87",x"c7"),
   593 => (x"c4",x"49",x"bf",x"ff"),
   594 => (x"ea",x"e2",x"c2",x"31"),
   595 => (x"87",x"ec",x"f6",x"59"),
   596 => (x"5c",x"5b",x"5e",x"0e"),
   597 => (x"c0",x"4a",x"71",x"0e"),
   598 => (x"02",x"9a",x"72",x"4b"),
   599 => (x"da",x"87",x"e0",x"c0"),
   600 => (x"69",x"9f",x"49",x"a2"),
   601 => (x"e2",x"e2",x"c2",x"4b"),
   602 => (x"87",x"cf",x"02",x"bf"),
   603 => (x"9f",x"49",x"a2",x"d4"),
   604 => (x"c0",x"4c",x"49",x"69"),
   605 => (x"d0",x"9c",x"ff",x"ff"),
   606 => (x"c0",x"87",x"c2",x"34"),
   607 => (x"73",x"b3",x"74",x"4c"),
   608 => (x"87",x"ee",x"fd",x"49"),
   609 => (x"0e",x"87",x"f3",x"f5"),
   610 => (x"5d",x"5c",x"5b",x"5e"),
   611 => (x"71",x"86",x"f4",x"0e"),
   612 => (x"72",x"7e",x"c0",x"4a"),
   613 => (x"87",x"d8",x"02",x"9a"),
   614 => (x"48",x"d6",x"da",x"c2"),
   615 => (x"da",x"c2",x"78",x"c0"),
   616 => (x"e7",x"c2",x"48",x"ce"),
   617 => (x"c2",x"78",x"bf",x"c7"),
   618 => (x"c2",x"48",x"d2",x"da"),
   619 => (x"78",x"bf",x"c3",x"e7"),
   620 => (x"48",x"f7",x"e2",x"c2"),
   621 => (x"e2",x"c2",x"50",x"c0"),
   622 => (x"c2",x"49",x"bf",x"e6"),
   623 => (x"4a",x"bf",x"d6",x"da"),
   624 => (x"c4",x"03",x"aa",x"71"),
   625 => (x"49",x"72",x"87",x"c9"),
   626 => (x"c0",x"05",x"99",x"cf"),
   627 => (x"ed",x"c0",x"87",x"e9"),
   628 => (x"da",x"c2",x"48",x"de"),
   629 => (x"c2",x"78",x"bf",x"ce"),
   630 => (x"c2",x"1e",x"da",x"da"),
   631 => (x"49",x"bf",x"ce",x"da"),
   632 => (x"48",x"ce",x"da",x"c2"),
   633 => (x"71",x"78",x"a1",x"c1"),
   634 => (x"c4",x"87",x"dd",x"e6"),
   635 => (x"da",x"ed",x"c0",x"86"),
   636 => (x"da",x"da",x"c2",x"48"),
   637 => (x"c0",x"87",x"cc",x"78"),
   638 => (x"48",x"bf",x"da",x"ed"),
   639 => (x"c0",x"80",x"e0",x"c0"),
   640 => (x"c2",x"58",x"de",x"ed"),
   641 => (x"48",x"bf",x"d6",x"da"),
   642 => (x"da",x"c2",x"80",x"c1"),
   643 => (x"5a",x"27",x"58",x"da"),
   644 => (x"bf",x"00",x"00",x"0b"),
   645 => (x"9d",x"4d",x"bf",x"97"),
   646 => (x"87",x"e3",x"c2",x"02"),
   647 => (x"02",x"ad",x"e5",x"c3"),
   648 => (x"c0",x"87",x"dc",x"c2"),
   649 => (x"4b",x"bf",x"da",x"ed"),
   650 => (x"11",x"49",x"a3",x"cb"),
   651 => (x"05",x"ac",x"cf",x"4c"),
   652 => (x"75",x"87",x"d2",x"c1"),
   653 => (x"c1",x"99",x"df",x"49"),
   654 => (x"c2",x"91",x"cd",x"89"),
   655 => (x"c1",x"81",x"ea",x"e2"),
   656 => (x"51",x"12",x"4a",x"a3"),
   657 => (x"12",x"4a",x"a3",x"c3"),
   658 => (x"4a",x"a3",x"c5",x"51"),
   659 => (x"a3",x"c7",x"51",x"12"),
   660 => (x"c9",x"51",x"12",x"4a"),
   661 => (x"51",x"12",x"4a",x"a3"),
   662 => (x"12",x"4a",x"a3",x"ce"),
   663 => (x"4a",x"a3",x"d0",x"51"),
   664 => (x"a3",x"d2",x"51",x"12"),
   665 => (x"d4",x"51",x"12",x"4a"),
   666 => (x"51",x"12",x"4a",x"a3"),
   667 => (x"12",x"4a",x"a3",x"d6"),
   668 => (x"4a",x"a3",x"d8",x"51"),
   669 => (x"a3",x"dc",x"51",x"12"),
   670 => (x"de",x"51",x"12",x"4a"),
   671 => (x"51",x"12",x"4a",x"a3"),
   672 => (x"fa",x"c0",x"7e",x"c1"),
   673 => (x"c8",x"49",x"74",x"87"),
   674 => (x"eb",x"c0",x"05",x"99"),
   675 => (x"d0",x"49",x"74",x"87"),
   676 => (x"87",x"d1",x"05",x"99"),
   677 => (x"c0",x"02",x"66",x"dc"),
   678 => (x"49",x"73",x"87",x"cb"),
   679 => (x"70",x"0f",x"66",x"dc"),
   680 => (x"d3",x"c0",x"02",x"98"),
   681 => (x"c0",x"05",x"6e",x"87"),
   682 => (x"e2",x"c2",x"87",x"c6"),
   683 => (x"50",x"c0",x"48",x"ea"),
   684 => (x"bf",x"da",x"ed",x"c0"),
   685 => (x"87",x"dd",x"c2",x"48"),
   686 => (x"48",x"f7",x"e2",x"c2"),
   687 => (x"c2",x"7e",x"50",x"c0"),
   688 => (x"49",x"bf",x"e6",x"e2"),
   689 => (x"bf",x"d6",x"da",x"c2"),
   690 => (x"04",x"aa",x"71",x"4a"),
   691 => (x"c2",x"87",x"f7",x"fb"),
   692 => (x"05",x"bf",x"c7",x"e7"),
   693 => (x"c2",x"87",x"c8",x"c0"),
   694 => (x"02",x"bf",x"e2",x"e2"),
   695 => (x"c2",x"87",x"f4",x"c1"),
   696 => (x"49",x"bf",x"d2",x"da"),
   697 => (x"c2",x"87",x"d9",x"f0"),
   698 => (x"c4",x"58",x"d6",x"da"),
   699 => (x"da",x"c2",x"48",x"a6"),
   700 => (x"c2",x"78",x"bf",x"d2"),
   701 => (x"02",x"bf",x"e2",x"e2"),
   702 => (x"c4",x"87",x"d8",x"c0"),
   703 => (x"ff",x"cf",x"49",x"66"),
   704 => (x"99",x"f8",x"ff",x"ff"),
   705 => (x"c5",x"c0",x"02",x"a9"),
   706 => (x"c0",x"4c",x"c0",x"87"),
   707 => (x"4c",x"c1",x"87",x"e1"),
   708 => (x"c4",x"87",x"dc",x"c0"),
   709 => (x"ff",x"cf",x"49",x"66"),
   710 => (x"02",x"a9",x"99",x"f8"),
   711 => (x"c8",x"87",x"c8",x"c0"),
   712 => (x"78",x"c0",x"48",x"a6"),
   713 => (x"c8",x"87",x"c5",x"c0"),
   714 => (x"78",x"c1",x"48",x"a6"),
   715 => (x"74",x"4c",x"66",x"c8"),
   716 => (x"de",x"c0",x"05",x"9c"),
   717 => (x"49",x"66",x"c4",x"87"),
   718 => (x"e2",x"c2",x"89",x"c2"),
   719 => (x"c2",x"91",x"bf",x"da"),
   720 => (x"48",x"bf",x"f3",x"e6"),
   721 => (x"da",x"c2",x"80",x"71"),
   722 => (x"da",x"c2",x"58",x"d2"),
   723 => (x"78",x"c0",x"48",x"d6"),
   724 => (x"c0",x"87",x"e3",x"f9"),
   725 => (x"ee",x"8e",x"f4",x"48"),
   726 => (x"00",x"00",x"87",x"de"),
   727 => (x"ff",x"ff",x"00",x"00"),
   728 => (x"0b",x"6a",x"ff",x"ff"),
   729 => (x"0b",x"73",x"00",x"00"),
   730 => (x"41",x"46",x"00",x"00"),
   731 => (x"20",x"32",x"33",x"54"),
   732 => (x"46",x"00",x"20",x"20"),
   733 => (x"36",x"31",x"54",x"41"),
   734 => (x"00",x"20",x"20",x"20"),
   735 => (x"48",x"d4",x"ff",x"1e"),
   736 => (x"68",x"78",x"ff",x"c3"),
   737 => (x"1e",x"4f",x"26",x"48"),
   738 => (x"c3",x"48",x"d4",x"ff"),
   739 => (x"d0",x"ff",x"78",x"ff"),
   740 => (x"78",x"e1",x"c0",x"48"),
   741 => (x"d4",x"48",x"d4",x"ff"),
   742 => (x"cb",x"e7",x"c2",x"78"),
   743 => (x"bf",x"d4",x"ff",x"48"),
   744 => (x"1e",x"4f",x"26",x"50"),
   745 => (x"c0",x"48",x"d0",x"ff"),
   746 => (x"4f",x"26",x"78",x"e0"),
   747 => (x"87",x"cc",x"ff",x"1e"),
   748 => (x"02",x"99",x"49",x"70"),
   749 => (x"fb",x"c0",x"87",x"c6"),
   750 => (x"87",x"f1",x"05",x"a9"),
   751 => (x"4f",x"26",x"48",x"71"),
   752 => (x"5c",x"5b",x"5e",x"0e"),
   753 => (x"c0",x"4b",x"71",x"0e"),
   754 => (x"87",x"f0",x"fe",x"4c"),
   755 => (x"02",x"99",x"49",x"70"),
   756 => (x"c0",x"87",x"f9",x"c0"),
   757 => (x"c0",x"02",x"a9",x"ec"),
   758 => (x"fb",x"c0",x"87",x"f2"),
   759 => (x"eb",x"c0",x"02",x"a9"),
   760 => (x"b7",x"66",x"cc",x"87"),
   761 => (x"87",x"c7",x"03",x"ac"),
   762 => (x"c2",x"02",x"66",x"d0"),
   763 => (x"71",x"53",x"71",x"87"),
   764 => (x"87",x"c2",x"02",x"99"),
   765 => (x"c3",x"fe",x"84",x"c1"),
   766 => (x"99",x"49",x"70",x"87"),
   767 => (x"c0",x"87",x"cd",x"02"),
   768 => (x"c7",x"02",x"a9",x"ec"),
   769 => (x"a9",x"fb",x"c0",x"87"),
   770 => (x"87",x"d5",x"ff",x"05"),
   771 => (x"c3",x"02",x"66",x"d0"),
   772 => (x"7b",x"97",x"c0",x"87"),
   773 => (x"05",x"a9",x"ec",x"c0"),
   774 => (x"4a",x"74",x"87",x"c4"),
   775 => (x"4a",x"74",x"87",x"c5"),
   776 => (x"72",x"8a",x"0a",x"c0"),
   777 => (x"26",x"87",x"c2",x"48"),
   778 => (x"26",x"4c",x"26",x"4d"),
   779 => (x"1e",x"4f",x"26",x"4b"),
   780 => (x"70",x"87",x"c9",x"fd"),
   781 => (x"aa",x"f0",x"c0",x"4a"),
   782 => (x"c0",x"87",x"c9",x"04"),
   783 => (x"c3",x"01",x"aa",x"f9"),
   784 => (x"8a",x"f0",x"c0",x"87"),
   785 => (x"04",x"aa",x"c1",x"c1"),
   786 => (x"da",x"c1",x"87",x"c9"),
   787 => (x"87",x"c3",x"01",x"aa"),
   788 => (x"72",x"8a",x"f7",x"c0"),
   789 => (x"0e",x"4f",x"26",x"48"),
   790 => (x"0e",x"5c",x"5b",x"5e"),
   791 => (x"d4",x"ff",x"4a",x"71"),
   792 => (x"c0",x"49",x"72",x"4b"),
   793 => (x"4c",x"70",x"87",x"e7"),
   794 => (x"87",x"c2",x"02",x"9c"),
   795 => (x"d0",x"ff",x"8c",x"c1"),
   796 => (x"c1",x"78",x"c5",x"48"),
   797 => (x"49",x"74",x"7b",x"d5"),
   798 => (x"de",x"c1",x"31",x"c6"),
   799 => (x"4a",x"bf",x"97",x"c5"),
   800 => (x"70",x"b0",x"71",x"48"),
   801 => (x"48",x"d0",x"ff",x"7b"),
   802 => (x"dc",x"fe",x"78",x"c4"),
   803 => (x"5b",x"5e",x"0e",x"87"),
   804 => (x"f8",x"0e",x"5d",x"5c"),
   805 => (x"c0",x"4c",x"71",x"86"),
   806 => (x"87",x"eb",x"fb",x"7e"),
   807 => (x"f4",x"c0",x"4b",x"c0"),
   808 => (x"49",x"bf",x"97",x"fa"),
   809 => (x"cf",x"04",x"a9",x"c0"),
   810 => (x"87",x"c0",x"fc",x"87"),
   811 => (x"f4",x"c0",x"83",x"c1"),
   812 => (x"49",x"bf",x"97",x"fa"),
   813 => (x"87",x"f1",x"06",x"ab"),
   814 => (x"97",x"fa",x"f4",x"c0"),
   815 => (x"87",x"cf",x"02",x"bf"),
   816 => (x"70",x"87",x"f9",x"fa"),
   817 => (x"c6",x"02",x"99",x"49"),
   818 => (x"a9",x"ec",x"c0",x"87"),
   819 => (x"c0",x"87",x"f1",x"05"),
   820 => (x"87",x"e8",x"fa",x"4b"),
   821 => (x"e3",x"fa",x"4d",x"70"),
   822 => (x"58",x"a6",x"c8",x"87"),
   823 => (x"70",x"87",x"dd",x"fa"),
   824 => (x"c8",x"83",x"c1",x"4a"),
   825 => (x"69",x"97",x"49",x"a4"),
   826 => (x"c7",x"02",x"ad",x"49"),
   827 => (x"ad",x"ff",x"c0",x"87"),
   828 => (x"87",x"e7",x"c0",x"05"),
   829 => (x"97",x"49",x"a4",x"c9"),
   830 => (x"66",x"c4",x"49",x"69"),
   831 => (x"87",x"c7",x"02",x"a9"),
   832 => (x"a8",x"ff",x"c0",x"48"),
   833 => (x"ca",x"87",x"d4",x"05"),
   834 => (x"69",x"97",x"49",x"a4"),
   835 => (x"c6",x"02",x"aa",x"49"),
   836 => (x"aa",x"ff",x"c0",x"87"),
   837 => (x"c1",x"87",x"c4",x"05"),
   838 => (x"c0",x"87",x"d0",x"7e"),
   839 => (x"c6",x"02",x"ad",x"ec"),
   840 => (x"ad",x"fb",x"c0",x"87"),
   841 => (x"c0",x"87",x"c4",x"05"),
   842 => (x"6e",x"7e",x"c1",x"4b"),
   843 => (x"87",x"e1",x"fe",x"02"),
   844 => (x"73",x"87",x"f0",x"f9"),
   845 => (x"fb",x"8e",x"f8",x"48"),
   846 => (x"0e",x"00",x"87",x"ed"),
   847 => (x"5d",x"5c",x"5b",x"5e"),
   848 => (x"71",x"86",x"f8",x"0e"),
   849 => (x"4b",x"d4",x"ff",x"4d"),
   850 => (x"e7",x"c2",x"1e",x"75"),
   851 => (x"e1",x"e8",x"49",x"d0"),
   852 => (x"70",x"86",x"c4",x"87"),
   853 => (x"ca",x"c4",x"02",x"98"),
   854 => (x"48",x"a6",x"c4",x"87"),
   855 => (x"bf",x"c7",x"de",x"c1"),
   856 => (x"fb",x"49",x"75",x"78"),
   857 => (x"d0",x"ff",x"87",x"f1"),
   858 => (x"c1",x"78",x"c5",x"48"),
   859 => (x"4a",x"c0",x"7b",x"d6"),
   860 => (x"11",x"49",x"a2",x"75"),
   861 => (x"cb",x"82",x"c1",x"7b"),
   862 => (x"f3",x"04",x"aa",x"b7"),
   863 => (x"c3",x"4a",x"cc",x"87"),
   864 => (x"82",x"c1",x"7b",x"ff"),
   865 => (x"aa",x"b7",x"e0",x"c0"),
   866 => (x"ff",x"87",x"f4",x"04"),
   867 => (x"78",x"c4",x"48",x"d0"),
   868 => (x"c5",x"7b",x"ff",x"c3"),
   869 => (x"7b",x"d3",x"c1",x"78"),
   870 => (x"78",x"c4",x"7b",x"c1"),
   871 => (x"b7",x"c0",x"48",x"66"),
   872 => (x"ee",x"c2",x"06",x"a8"),
   873 => (x"d8",x"e7",x"c2",x"87"),
   874 => (x"66",x"c4",x"4c",x"bf"),
   875 => (x"c8",x"88",x"74",x"48"),
   876 => (x"9c",x"74",x"58",x"a6"),
   877 => (x"87",x"f7",x"c1",x"02"),
   878 => (x"7e",x"da",x"da",x"c2"),
   879 => (x"8c",x"4d",x"c0",x"c8"),
   880 => (x"03",x"ac",x"b7",x"c0"),
   881 => (x"c0",x"c8",x"87",x"c6"),
   882 => (x"4c",x"c0",x"4d",x"a4"),
   883 => (x"97",x"cb",x"e7",x"c2"),
   884 => (x"99",x"d0",x"49",x"bf"),
   885 => (x"c0",x"87",x"d0",x"02"),
   886 => (x"d0",x"e7",x"c2",x"1e"),
   887 => (x"87",x"c4",x"eb",x"49"),
   888 => (x"4a",x"70",x"86",x"c4"),
   889 => (x"c2",x"87",x"ed",x"c0"),
   890 => (x"c2",x"1e",x"da",x"da"),
   891 => (x"ea",x"49",x"d0",x"e7"),
   892 => (x"86",x"c4",x"87",x"f2"),
   893 => (x"d0",x"ff",x"4a",x"70"),
   894 => (x"78",x"c5",x"c8",x"48"),
   895 => (x"6e",x"7b",x"d4",x"c1"),
   896 => (x"6e",x"7b",x"bf",x"97"),
   897 => (x"70",x"80",x"c1",x"48"),
   898 => (x"05",x"8d",x"c1",x"7e"),
   899 => (x"ff",x"87",x"f0",x"ff"),
   900 => (x"78",x"c4",x"48",x"d0"),
   901 => (x"c5",x"05",x"9a",x"72"),
   902 => (x"c1",x"48",x"c0",x"87"),
   903 => (x"1e",x"c1",x"87",x"c7"),
   904 => (x"49",x"d0",x"e7",x"c2"),
   905 => (x"c4",x"87",x"e3",x"e8"),
   906 => (x"05",x"9c",x"74",x"86"),
   907 => (x"c4",x"87",x"c9",x"fe"),
   908 => (x"b7",x"c0",x"48",x"66"),
   909 => (x"87",x"d1",x"06",x"a8"),
   910 => (x"48",x"d0",x"e7",x"c2"),
   911 => (x"80",x"d0",x"78",x"c0"),
   912 => (x"80",x"f4",x"78",x"c0"),
   913 => (x"bf",x"dc",x"e7",x"c2"),
   914 => (x"48",x"66",x"c4",x"78"),
   915 => (x"01",x"a8",x"b7",x"c0"),
   916 => (x"ff",x"87",x"d2",x"fd"),
   917 => (x"78",x"c5",x"48",x"d0"),
   918 => (x"c0",x"7b",x"d3",x"c1"),
   919 => (x"c1",x"78",x"c4",x"7b"),
   920 => (x"c0",x"87",x"c2",x"48"),
   921 => (x"26",x"8e",x"f8",x"48"),
   922 => (x"26",x"4c",x"26",x"4d"),
   923 => (x"0e",x"4f",x"26",x"4b"),
   924 => (x"5d",x"5c",x"5b",x"5e"),
   925 => (x"4b",x"71",x"1e",x"0e"),
   926 => (x"ab",x"4d",x"4c",x"c0"),
   927 => (x"87",x"e8",x"c0",x"04"),
   928 => (x"1e",x"cd",x"f2",x"c0"),
   929 => (x"c4",x"02",x"9d",x"75"),
   930 => (x"c2",x"4a",x"c0",x"87"),
   931 => (x"72",x"4a",x"c1",x"87"),
   932 => (x"87",x"f3",x"eb",x"49"),
   933 => (x"7e",x"70",x"86",x"c4"),
   934 => (x"05",x"6e",x"84",x"c1"),
   935 => (x"4c",x"73",x"87",x"c2"),
   936 => (x"ac",x"73",x"85",x"c1"),
   937 => (x"87",x"d8",x"ff",x"06"),
   938 => (x"fe",x"26",x"48",x"6e"),
   939 => (x"71",x"1e",x"87",x"f9"),
   940 => (x"05",x"66",x"c4",x"4a"),
   941 => (x"49",x"72",x"87",x"c5"),
   942 => (x"26",x"87",x"c0",x"fa"),
   943 => (x"5b",x"5e",x"0e",x"4f"),
   944 => (x"1e",x"0e",x"5d",x"5c"),
   945 => (x"de",x"49",x"4c",x"71"),
   946 => (x"f8",x"e7",x"c2",x"91"),
   947 => (x"97",x"85",x"71",x"4d"),
   948 => (x"dc",x"c1",x"02",x"6d"),
   949 => (x"e4",x"e7",x"c2",x"87"),
   950 => (x"81",x"74",x"49",x"bf"),
   951 => (x"87",x"cf",x"fe",x"71"),
   952 => (x"98",x"48",x"7e",x"70"),
   953 => (x"87",x"f2",x"c0",x"02"),
   954 => (x"4b",x"ec",x"e7",x"c2"),
   955 => (x"49",x"cb",x"4a",x"70"),
   956 => (x"87",x"f3",x"c6",x"ff"),
   957 => (x"93",x"cb",x"4b",x"74"),
   958 => (x"83",x"d9",x"de",x"c1"),
   959 => (x"fc",x"c0",x"83",x"c4"),
   960 => (x"49",x"74",x"7b",x"f5"),
   961 => (x"87",x"ce",x"cd",x"c1"),
   962 => (x"de",x"c1",x"7b",x"75"),
   963 => (x"49",x"bf",x"97",x"c6"),
   964 => (x"ec",x"e7",x"c2",x"1e"),
   965 => (x"87",x"d6",x"fe",x"49"),
   966 => (x"49",x"74",x"86",x"c4"),
   967 => (x"87",x"f6",x"cc",x"c1"),
   968 => (x"ce",x"c1",x"49",x"c0"),
   969 => (x"e7",x"c2",x"87",x"d5"),
   970 => (x"78",x"c0",x"48",x"cc"),
   971 => (x"f9",x"dd",x"49",x"c1"),
   972 => (x"f2",x"fc",x"26",x"87"),
   973 => (x"61",x"6f",x"4c",x"87"),
   974 => (x"67",x"6e",x"69",x"64"),
   975 => (x"00",x"2e",x"2e",x"2e"),
   976 => (x"71",x"1e",x"73",x"1e"),
   977 => (x"e7",x"c2",x"49",x"4a"),
   978 => (x"71",x"81",x"bf",x"e4"),
   979 => (x"70",x"87",x"e0",x"fc"),
   980 => (x"c4",x"02",x"9b",x"4b"),
   981 => (x"f7",x"e7",x"49",x"87"),
   982 => (x"e4",x"e7",x"c2",x"87"),
   983 => (x"c1",x"78",x"c0",x"48"),
   984 => (x"87",x"c6",x"dd",x"49"),
   985 => (x"1e",x"87",x"c4",x"fc"),
   986 => (x"cd",x"c1",x"49",x"c0"),
   987 => (x"4f",x"26",x"87",x"cd"),
   988 => (x"49",x"4a",x"71",x"1e"),
   989 => (x"de",x"c1",x"91",x"cb"),
   990 => (x"81",x"c8",x"81",x"d9"),
   991 => (x"e7",x"c2",x"48",x"11"),
   992 => (x"e7",x"c2",x"58",x"d0"),
   993 => (x"78",x"c0",x"48",x"e4"),
   994 => (x"dd",x"dc",x"49",x"c1"),
   995 => (x"1e",x"4f",x"26",x"87"),
   996 => (x"d2",x"02",x"99",x"71"),
   997 => (x"ee",x"df",x"c1",x"87"),
   998 => (x"f7",x"50",x"c0",x"48"),
   999 => (x"f0",x"fd",x"c0",x"80"),
  1000 => (x"d2",x"de",x"c1",x"40"),
  1001 => (x"c1",x"87",x"ce",x"78"),
  1002 => (x"c1",x"48",x"ea",x"df"),
  1003 => (x"fc",x"78",x"cb",x"de"),
  1004 => (x"e7",x"fd",x"c0",x"80"),
  1005 => (x"0e",x"4f",x"26",x"78"),
  1006 => (x"5d",x"5c",x"5b",x"5e"),
  1007 => (x"c2",x"86",x"f4",x"0e"),
  1008 => (x"c0",x"4d",x"da",x"da"),
  1009 => (x"48",x"a6",x"c4",x"4c"),
  1010 => (x"e7",x"c2",x"78",x"c0"),
  1011 => (x"c0",x"48",x"bf",x"e4"),
  1012 => (x"c0",x"c1",x"06",x"a8"),
  1013 => (x"da",x"da",x"c2",x"87"),
  1014 => (x"c0",x"02",x"98",x"48"),
  1015 => (x"f2",x"c0",x"87",x"f7"),
  1016 => (x"66",x"c8",x"1e",x"cd"),
  1017 => (x"c4",x"87",x"c7",x"02"),
  1018 => (x"78",x"c0",x"48",x"a6"),
  1019 => (x"a6",x"c4",x"87",x"c5"),
  1020 => (x"c4",x"78",x"c1",x"48"),
  1021 => (x"ce",x"e6",x"49",x"66"),
  1022 => (x"70",x"86",x"c4",x"87"),
  1023 => (x"c4",x"84",x"c1",x"4d"),
  1024 => (x"80",x"c1",x"48",x"66"),
  1025 => (x"c2",x"58",x"a6",x"c8"),
  1026 => (x"ac",x"bf",x"e4",x"e7"),
  1027 => (x"75",x"87",x"c6",x"03"),
  1028 => (x"c9",x"ff",x"05",x"9d"),
  1029 => (x"75",x"4c",x"c0",x"87"),
  1030 => (x"dc",x"c3",x"02",x"9d"),
  1031 => (x"cd",x"f2",x"c0",x"87"),
  1032 => (x"02",x"66",x"c8",x"1e"),
  1033 => (x"a6",x"cc",x"87",x"c7"),
  1034 => (x"c5",x"78",x"c0",x"48"),
  1035 => (x"48",x"a6",x"cc",x"87"),
  1036 => (x"66",x"cc",x"78",x"c1"),
  1037 => (x"87",x"cf",x"e5",x"49"),
  1038 => (x"7e",x"70",x"86",x"c4"),
  1039 => (x"c2",x"02",x"98",x"48"),
  1040 => (x"cb",x"49",x"87",x"e4"),
  1041 => (x"49",x"69",x"97",x"81"),
  1042 => (x"c1",x"02",x"99",x"d0"),
  1043 => (x"49",x"74",x"87",x"d4"),
  1044 => (x"de",x"c1",x"91",x"cb"),
  1045 => (x"fd",x"c0",x"81",x"d9"),
  1046 => (x"81",x"c8",x"79",x"c0"),
  1047 => (x"74",x"51",x"ff",x"c3"),
  1048 => (x"c2",x"91",x"de",x"49"),
  1049 => (x"71",x"4d",x"f8",x"e7"),
  1050 => (x"97",x"c1",x"c2",x"85"),
  1051 => (x"49",x"a5",x"c1",x"7d"),
  1052 => (x"c2",x"51",x"e0",x"c0"),
  1053 => (x"bf",x"97",x"ea",x"e2"),
  1054 => (x"c1",x"87",x"d2",x"02"),
  1055 => (x"4b",x"a5",x"c2",x"84"),
  1056 => (x"4a",x"ea",x"e2",x"c2"),
  1057 => (x"c0",x"ff",x"49",x"db"),
  1058 => (x"d9",x"c1",x"87",x"dd"),
  1059 => (x"49",x"a5",x"cd",x"87"),
  1060 => (x"84",x"c1",x"51",x"c0"),
  1061 => (x"6e",x"4b",x"a5",x"c2"),
  1062 => (x"ff",x"49",x"cb",x"4a"),
  1063 => (x"c1",x"87",x"c8",x"c0"),
  1064 => (x"49",x"74",x"87",x"c4"),
  1065 => (x"de",x"c1",x"91",x"cb"),
  1066 => (x"fa",x"c0",x"81",x"d9"),
  1067 => (x"e2",x"c2",x"79",x"fd"),
  1068 => (x"02",x"bf",x"97",x"ea"),
  1069 => (x"49",x"74",x"87",x"d8"),
  1070 => (x"84",x"c1",x"91",x"de"),
  1071 => (x"4b",x"f8",x"e7",x"c2"),
  1072 => (x"e2",x"c2",x"83",x"71"),
  1073 => (x"49",x"dd",x"4a",x"ea"),
  1074 => (x"87",x"db",x"ff",x"fe"),
  1075 => (x"4b",x"74",x"87",x"d8"),
  1076 => (x"e7",x"c2",x"93",x"de"),
  1077 => (x"a3",x"cb",x"83",x"f8"),
  1078 => (x"c1",x"51",x"c0",x"49"),
  1079 => (x"4a",x"6e",x"73",x"84"),
  1080 => (x"ff",x"fe",x"49",x"cb"),
  1081 => (x"66",x"c4",x"87",x"c1"),
  1082 => (x"c8",x"80",x"c1",x"48"),
  1083 => (x"ac",x"c7",x"58",x"a6"),
  1084 => (x"87",x"c5",x"c0",x"03"),
  1085 => (x"e4",x"fc",x"05",x"6e"),
  1086 => (x"f4",x"48",x"74",x"87"),
  1087 => (x"87",x"e7",x"f5",x"8e"),
  1088 => (x"71",x"1e",x"73",x"1e"),
  1089 => (x"91",x"cb",x"49",x"4b"),
  1090 => (x"81",x"d9",x"de",x"c1"),
  1091 => (x"c1",x"4a",x"a1",x"c8"),
  1092 => (x"12",x"48",x"c5",x"de"),
  1093 => (x"4a",x"a1",x"c9",x"50"),
  1094 => (x"48",x"fa",x"f4",x"c0"),
  1095 => (x"81",x"ca",x"50",x"12"),
  1096 => (x"48",x"c6",x"de",x"c1"),
  1097 => (x"de",x"c1",x"50",x"11"),
  1098 => (x"49",x"bf",x"97",x"c6"),
  1099 => (x"f5",x"49",x"c0",x"1e"),
  1100 => (x"e7",x"c2",x"87",x"fc"),
  1101 => (x"78",x"de",x"48",x"cc"),
  1102 => (x"ed",x"d5",x"49",x"c1"),
  1103 => (x"ea",x"f4",x"26",x"87"),
  1104 => (x"5b",x"5e",x"0e",x"87"),
  1105 => (x"f4",x"0e",x"5d",x"5c"),
  1106 => (x"49",x"4d",x"71",x"86"),
  1107 => (x"de",x"c1",x"91",x"cb"),
  1108 => (x"a1",x"c8",x"81",x"d9"),
  1109 => (x"7e",x"a1",x"ca",x"4a"),
  1110 => (x"c2",x"48",x"a6",x"c4"),
  1111 => (x"78",x"bf",x"fa",x"eb"),
  1112 => (x"4b",x"bf",x"97",x"6e"),
  1113 => (x"73",x"4c",x"66",x"c4"),
  1114 => (x"cc",x"48",x"12",x"2c"),
  1115 => (x"9c",x"70",x"58",x"a6"),
  1116 => (x"81",x"c9",x"84",x"c1"),
  1117 => (x"b7",x"49",x"69",x"97"),
  1118 => (x"87",x"c2",x"04",x"ac"),
  1119 => (x"97",x"6e",x"4c",x"c0"),
  1120 => (x"66",x"c8",x"4a",x"bf"),
  1121 => (x"ff",x"31",x"72",x"49"),
  1122 => (x"99",x"66",x"c4",x"b9"),
  1123 => (x"30",x"72",x"48",x"74"),
  1124 => (x"71",x"48",x"4a",x"70"),
  1125 => (x"fe",x"eb",x"c2",x"b0"),
  1126 => (x"f9",x"f0",x"c0",x"58"),
  1127 => (x"d4",x"49",x"c0",x"87"),
  1128 => (x"49",x"75",x"87",x"c8"),
  1129 => (x"87",x"ee",x"c2",x"c1"),
  1130 => (x"fa",x"f2",x"8e",x"f4"),
  1131 => (x"1e",x"73",x"1e",x"87"),
  1132 => (x"fe",x"49",x"4b",x"71"),
  1133 => (x"49",x"73",x"87",x"cb"),
  1134 => (x"f2",x"87",x"c6",x"fe"),
  1135 => (x"73",x"1e",x"87",x"ed"),
  1136 => (x"c6",x"4b",x"71",x"1e"),
  1137 => (x"db",x"02",x"4a",x"a3"),
  1138 => (x"02",x"8a",x"c1",x"87"),
  1139 => (x"02",x"8a",x"87",x"d6"),
  1140 => (x"8a",x"87",x"da",x"c1"),
  1141 => (x"87",x"fc",x"c0",x"02"),
  1142 => (x"e1",x"c0",x"02",x"8a"),
  1143 => (x"cb",x"02",x"8a",x"87"),
  1144 => (x"87",x"db",x"c1",x"87"),
  1145 => (x"c7",x"f6",x"49",x"c7"),
  1146 => (x"87",x"de",x"c1",x"87"),
  1147 => (x"bf",x"e4",x"e7",x"c2"),
  1148 => (x"87",x"cb",x"c1",x"02"),
  1149 => (x"c2",x"88",x"c1",x"48"),
  1150 => (x"c1",x"58",x"e8",x"e7"),
  1151 => (x"e7",x"c2",x"87",x"c1"),
  1152 => (x"c0",x"02",x"bf",x"e8"),
  1153 => (x"e7",x"c2",x"87",x"f9"),
  1154 => (x"c1",x"48",x"bf",x"e4"),
  1155 => (x"e8",x"e7",x"c2",x"80"),
  1156 => (x"87",x"eb",x"c0",x"58"),
  1157 => (x"bf",x"e4",x"e7",x"c2"),
  1158 => (x"c2",x"89",x"c6",x"49"),
  1159 => (x"c0",x"59",x"e8",x"e7"),
  1160 => (x"da",x"03",x"a9",x"b7"),
  1161 => (x"e4",x"e7",x"c2",x"87"),
  1162 => (x"d2",x"78",x"c0",x"48"),
  1163 => (x"e8",x"e7",x"c2",x"87"),
  1164 => (x"87",x"cb",x"02",x"bf"),
  1165 => (x"bf",x"e4",x"e7",x"c2"),
  1166 => (x"c2",x"80",x"c6",x"48"),
  1167 => (x"c0",x"58",x"e8",x"e7"),
  1168 => (x"87",x"e6",x"d1",x"49"),
  1169 => (x"c0",x"c1",x"49",x"73"),
  1170 => (x"de",x"f0",x"87",x"cc"),
  1171 => (x"5b",x"5e",x"0e",x"87"),
  1172 => (x"ff",x"0e",x"5d",x"5c"),
  1173 => (x"a6",x"dc",x"86",x"d4"),
  1174 => (x"48",x"a6",x"c8",x"59"),
  1175 => (x"80",x"c4",x"78",x"c0"),
  1176 => (x"78",x"66",x"c0",x"c1"),
  1177 => (x"78",x"c1",x"80",x"c4"),
  1178 => (x"78",x"c1",x"80",x"c4"),
  1179 => (x"48",x"e8",x"e7",x"c2"),
  1180 => (x"e7",x"c2",x"78",x"c1"),
  1181 => (x"de",x"48",x"bf",x"cc"),
  1182 => (x"87",x"c9",x"05",x"a8"),
  1183 => (x"cc",x"87",x"f8",x"f4"),
  1184 => (x"e4",x"cf",x"58",x"a6"),
  1185 => (x"87",x"ff",x"e3",x"87"),
  1186 => (x"e3",x"87",x"e1",x"e4"),
  1187 => (x"4c",x"70",x"87",x"ee"),
  1188 => (x"02",x"ac",x"fb",x"c0"),
  1189 => (x"d8",x"87",x"fb",x"c1"),
  1190 => (x"ed",x"c1",x"05",x"66"),
  1191 => (x"66",x"fc",x"c0",x"87"),
  1192 => (x"6a",x"82",x"c4",x"4a"),
  1193 => (x"c1",x"1e",x"72",x"7e"),
  1194 => (x"c4",x"48",x"de",x"da"),
  1195 => (x"a1",x"c8",x"49",x"66"),
  1196 => (x"71",x"41",x"20",x"4a"),
  1197 => (x"87",x"f9",x"05",x"aa"),
  1198 => (x"4a",x"26",x"51",x"10"),
  1199 => (x"48",x"66",x"fc",x"c0"),
  1200 => (x"78",x"c0",x"c4",x"c1"),
  1201 => (x"81",x"c7",x"49",x"6a"),
  1202 => (x"fc",x"c0",x"51",x"74"),
  1203 => (x"81",x"c8",x"49",x"66"),
  1204 => (x"fc",x"c0",x"51",x"c1"),
  1205 => (x"81",x"c9",x"49",x"66"),
  1206 => (x"fc",x"c0",x"51",x"c0"),
  1207 => (x"81",x"ca",x"49",x"66"),
  1208 => (x"1e",x"c1",x"51",x"c0"),
  1209 => (x"49",x"6a",x"1e",x"d8"),
  1210 => (x"d3",x"e3",x"81",x"c8"),
  1211 => (x"c1",x"86",x"c8",x"87"),
  1212 => (x"c0",x"48",x"66",x"c0"),
  1213 => (x"87",x"c7",x"01",x"a8"),
  1214 => (x"c1",x"48",x"a6",x"c8"),
  1215 => (x"c1",x"87",x"ce",x"78"),
  1216 => (x"c1",x"48",x"66",x"c0"),
  1217 => (x"58",x"a6",x"d0",x"88"),
  1218 => (x"df",x"e2",x"87",x"c3"),
  1219 => (x"48",x"a6",x"d0",x"87"),
  1220 => (x"9c",x"74",x"78",x"c2"),
  1221 => (x"87",x"cd",x"cd",x"02"),
  1222 => (x"c1",x"48",x"66",x"c8"),
  1223 => (x"03",x"a8",x"66",x"c4"),
  1224 => (x"dc",x"87",x"c2",x"cd"),
  1225 => (x"78",x"c0",x"48",x"a6"),
  1226 => (x"78",x"c0",x"80",x"e8"),
  1227 => (x"70",x"87",x"cd",x"e1"),
  1228 => (x"ac",x"d0",x"c1",x"4c"),
  1229 => (x"87",x"d5",x"c2",x"05"),
  1230 => (x"e3",x"7e",x"66",x"c4"),
  1231 => (x"a6",x"c8",x"87",x"f1"),
  1232 => (x"87",x"f8",x"e0",x"58"),
  1233 => (x"ec",x"c0",x"4c",x"70"),
  1234 => (x"eb",x"c1",x"05",x"ac"),
  1235 => (x"49",x"66",x"c8",x"87"),
  1236 => (x"fc",x"c0",x"91",x"cb"),
  1237 => (x"a1",x"c4",x"81",x"66"),
  1238 => (x"c8",x"4d",x"6a",x"4a"),
  1239 => (x"66",x"c4",x"4a",x"a1"),
  1240 => (x"f0",x"fd",x"c0",x"52"),
  1241 => (x"87",x"d4",x"e0",x"79"),
  1242 => (x"02",x"9c",x"4c",x"70"),
  1243 => (x"fb",x"c0",x"87",x"d8"),
  1244 => (x"87",x"d2",x"02",x"ac"),
  1245 => (x"c3",x"e0",x"55",x"74"),
  1246 => (x"9c",x"4c",x"70",x"87"),
  1247 => (x"c0",x"87",x"c7",x"02"),
  1248 => (x"ff",x"05",x"ac",x"fb"),
  1249 => (x"e0",x"c0",x"87",x"ee"),
  1250 => (x"55",x"c1",x"c2",x"55"),
  1251 => (x"d8",x"7d",x"97",x"c0"),
  1252 => (x"a8",x"6e",x"48",x"66"),
  1253 => (x"c8",x"87",x"db",x"05"),
  1254 => (x"66",x"cc",x"48",x"66"),
  1255 => (x"87",x"ca",x"04",x"a8"),
  1256 => (x"c1",x"48",x"66",x"c8"),
  1257 => (x"58",x"a6",x"cc",x"80"),
  1258 => (x"66",x"cc",x"87",x"c8"),
  1259 => (x"d0",x"88",x"c1",x"48"),
  1260 => (x"df",x"ff",x"58",x"a6"),
  1261 => (x"4c",x"70",x"87",x"c6"),
  1262 => (x"05",x"ac",x"d0",x"c1"),
  1263 => (x"66",x"d4",x"87",x"c8"),
  1264 => (x"d8",x"80",x"c1",x"48"),
  1265 => (x"d0",x"c1",x"58",x"a6"),
  1266 => (x"eb",x"fd",x"02",x"ac"),
  1267 => (x"48",x"66",x"c4",x"87"),
  1268 => (x"05",x"a8",x"66",x"d8"),
  1269 => (x"c0",x"87",x"e0",x"c9"),
  1270 => (x"c0",x"48",x"a6",x"e0"),
  1271 => (x"c0",x"48",x"74",x"78"),
  1272 => (x"7e",x"70",x"88",x"fb"),
  1273 => (x"c9",x"02",x"98",x"48"),
  1274 => (x"cb",x"48",x"87",x"e2"),
  1275 => (x"48",x"7e",x"70",x"88"),
  1276 => (x"cd",x"c1",x"02",x"98"),
  1277 => (x"88",x"c9",x"48",x"87"),
  1278 => (x"98",x"48",x"7e",x"70"),
  1279 => (x"87",x"fe",x"c3",x"02"),
  1280 => (x"70",x"88",x"c4",x"48"),
  1281 => (x"02",x"98",x"48",x"7e"),
  1282 => (x"c1",x"48",x"87",x"ce"),
  1283 => (x"48",x"7e",x"70",x"88"),
  1284 => (x"e9",x"c3",x"02",x"98"),
  1285 => (x"87",x"d6",x"c8",x"87"),
  1286 => (x"c0",x"48",x"a6",x"dc"),
  1287 => (x"dd",x"ff",x"78",x"f0"),
  1288 => (x"4c",x"70",x"87",x"da"),
  1289 => (x"02",x"ac",x"ec",x"c0"),
  1290 => (x"c0",x"87",x"c4",x"c0"),
  1291 => (x"c0",x"5c",x"a6",x"e0"),
  1292 => (x"cd",x"02",x"ac",x"ec"),
  1293 => (x"c3",x"dd",x"ff",x"87"),
  1294 => (x"c0",x"4c",x"70",x"87"),
  1295 => (x"ff",x"05",x"ac",x"ec"),
  1296 => (x"ec",x"c0",x"87",x"f3"),
  1297 => (x"c4",x"c0",x"02",x"ac"),
  1298 => (x"ef",x"dc",x"ff",x"87"),
  1299 => (x"ca",x"1e",x"c0",x"87"),
  1300 => (x"49",x"66",x"d0",x"1e"),
  1301 => (x"c4",x"c1",x"91",x"cb"),
  1302 => (x"80",x"71",x"48",x"66"),
  1303 => (x"c8",x"58",x"a6",x"cc"),
  1304 => (x"80",x"c4",x"48",x"66"),
  1305 => (x"cc",x"58",x"a6",x"d0"),
  1306 => (x"ff",x"49",x"bf",x"66"),
  1307 => (x"c1",x"87",x"d1",x"dd"),
  1308 => (x"d4",x"1e",x"de",x"1e"),
  1309 => (x"ff",x"49",x"bf",x"66"),
  1310 => (x"d0",x"87",x"c5",x"dd"),
  1311 => (x"48",x"49",x"70",x"86"),
  1312 => (x"c0",x"88",x"08",x"c0"),
  1313 => (x"c0",x"58",x"a6",x"e8"),
  1314 => (x"ee",x"c0",x"06",x"a8"),
  1315 => (x"66",x"e4",x"c0",x"87"),
  1316 => (x"03",x"a8",x"dd",x"48"),
  1317 => (x"c4",x"87",x"e4",x"c0"),
  1318 => (x"c0",x"49",x"bf",x"66"),
  1319 => (x"c0",x"81",x"66",x"e4"),
  1320 => (x"e4",x"c0",x"51",x"e0"),
  1321 => (x"81",x"c1",x"49",x"66"),
  1322 => (x"81",x"bf",x"66",x"c4"),
  1323 => (x"c0",x"51",x"c1",x"c2"),
  1324 => (x"c2",x"49",x"66",x"e4"),
  1325 => (x"bf",x"66",x"c4",x"81"),
  1326 => (x"6e",x"51",x"c0",x"81"),
  1327 => (x"c0",x"c4",x"c1",x"48"),
  1328 => (x"c8",x"49",x"6e",x"78"),
  1329 => (x"51",x"66",x"d0",x"81"),
  1330 => (x"81",x"c9",x"49",x"6e"),
  1331 => (x"6e",x"51",x"66",x"d4"),
  1332 => (x"dc",x"81",x"ca",x"49"),
  1333 => (x"66",x"d0",x"51",x"66"),
  1334 => (x"d4",x"80",x"c1",x"48"),
  1335 => (x"66",x"c8",x"58",x"a6"),
  1336 => (x"a8",x"66",x"cc",x"48"),
  1337 => (x"87",x"cb",x"c0",x"04"),
  1338 => (x"c1",x"48",x"66",x"c8"),
  1339 => (x"58",x"a6",x"cc",x"80"),
  1340 => (x"cc",x"87",x"d9",x"c5"),
  1341 => (x"88",x"c1",x"48",x"66"),
  1342 => (x"c5",x"58",x"a6",x"d0"),
  1343 => (x"dc",x"ff",x"87",x"ce"),
  1344 => (x"e8",x"c0",x"87",x"ed"),
  1345 => (x"dc",x"ff",x"58",x"a6"),
  1346 => (x"e0",x"c0",x"87",x"e5"),
  1347 => (x"ec",x"c0",x"58",x"a6"),
  1348 => (x"ca",x"c0",x"05",x"a8"),
  1349 => (x"48",x"a6",x"dc",x"87"),
  1350 => (x"78",x"66",x"e4",x"c0"),
  1351 => (x"ff",x"87",x"c4",x"c0"),
  1352 => (x"c8",x"87",x"d9",x"d9"),
  1353 => (x"91",x"cb",x"49",x"66"),
  1354 => (x"48",x"66",x"fc",x"c0"),
  1355 => (x"7e",x"70",x"80",x"71"),
  1356 => (x"6e",x"82",x"c8",x"4a"),
  1357 => (x"c0",x"81",x"ca",x"49"),
  1358 => (x"dc",x"51",x"66",x"e4"),
  1359 => (x"81",x"c1",x"49",x"66"),
  1360 => (x"89",x"66",x"e4",x"c0"),
  1361 => (x"30",x"71",x"48",x"c1"),
  1362 => (x"89",x"c1",x"49",x"70"),
  1363 => (x"c2",x"7a",x"97",x"71"),
  1364 => (x"49",x"bf",x"fa",x"eb"),
  1365 => (x"29",x"66",x"e4",x"c0"),
  1366 => (x"48",x"4a",x"6a",x"97"),
  1367 => (x"ec",x"c0",x"98",x"71"),
  1368 => (x"49",x"6e",x"58",x"a6"),
  1369 => (x"4d",x"69",x"81",x"c4"),
  1370 => (x"c4",x"48",x"66",x"d8"),
  1371 => (x"c0",x"02",x"a8",x"66"),
  1372 => (x"a6",x"c4",x"87",x"c8"),
  1373 => (x"c0",x"78",x"c0",x"48"),
  1374 => (x"a6",x"c4",x"87",x"c5"),
  1375 => (x"c4",x"78",x"c1",x"48"),
  1376 => (x"e0",x"c0",x"1e",x"66"),
  1377 => (x"ff",x"49",x"75",x"1e"),
  1378 => (x"c8",x"87",x"f5",x"d8"),
  1379 => (x"c0",x"4c",x"70",x"86"),
  1380 => (x"c1",x"06",x"ac",x"b7"),
  1381 => (x"85",x"74",x"87",x"d4"),
  1382 => (x"74",x"49",x"e0",x"c0"),
  1383 => (x"c1",x"4b",x"75",x"89"),
  1384 => (x"71",x"4a",x"e7",x"da"),
  1385 => (x"87",x"ff",x"eb",x"fe"),
  1386 => (x"e0",x"c0",x"85",x"c2"),
  1387 => (x"80",x"c1",x"48",x"66"),
  1388 => (x"58",x"a6",x"e4",x"c0"),
  1389 => (x"49",x"66",x"e8",x"c0"),
  1390 => (x"a9",x"70",x"81",x"c1"),
  1391 => (x"87",x"c8",x"c0",x"02"),
  1392 => (x"c0",x"48",x"a6",x"c4"),
  1393 => (x"87",x"c5",x"c0",x"78"),
  1394 => (x"c1",x"48",x"a6",x"c4"),
  1395 => (x"1e",x"66",x"c4",x"78"),
  1396 => (x"c0",x"49",x"a4",x"c2"),
  1397 => (x"88",x"71",x"48",x"e0"),
  1398 => (x"75",x"1e",x"49",x"70"),
  1399 => (x"df",x"d7",x"ff",x"49"),
  1400 => (x"c0",x"86",x"c8",x"87"),
  1401 => (x"ff",x"01",x"a8",x"b7"),
  1402 => (x"e0",x"c0",x"87",x"c0"),
  1403 => (x"d1",x"c0",x"02",x"66"),
  1404 => (x"c9",x"49",x"6e",x"87"),
  1405 => (x"66",x"e0",x"c0",x"81"),
  1406 => (x"c1",x"48",x"6e",x"51"),
  1407 => (x"c0",x"78",x"c1",x"c5"),
  1408 => (x"49",x"6e",x"87",x"cc"),
  1409 => (x"51",x"c2",x"81",x"c9"),
  1410 => (x"c6",x"c1",x"48",x"6e"),
  1411 => (x"66",x"c8",x"78",x"ed"),
  1412 => (x"a8",x"66",x"cc",x"48"),
  1413 => (x"87",x"cb",x"c0",x"04"),
  1414 => (x"c1",x"48",x"66",x"c8"),
  1415 => (x"58",x"a6",x"cc",x"80"),
  1416 => (x"cc",x"87",x"e9",x"c0"),
  1417 => (x"88",x"c1",x"48",x"66"),
  1418 => (x"c0",x"58",x"a6",x"d0"),
  1419 => (x"d5",x"ff",x"87",x"de"),
  1420 => (x"4c",x"70",x"87",x"fa"),
  1421 => (x"c1",x"87",x"d5",x"c0"),
  1422 => (x"c0",x"05",x"ac",x"c6"),
  1423 => (x"66",x"d0",x"87",x"c8"),
  1424 => (x"d4",x"80",x"c1",x"48"),
  1425 => (x"d5",x"ff",x"58",x"a6"),
  1426 => (x"4c",x"70",x"87",x"e2"),
  1427 => (x"c1",x"48",x"66",x"d4"),
  1428 => (x"58",x"a6",x"d8",x"80"),
  1429 => (x"c0",x"02",x"9c",x"74"),
  1430 => (x"66",x"c8",x"87",x"cb"),
  1431 => (x"66",x"c4",x"c1",x"48"),
  1432 => (x"fe",x"f2",x"04",x"a8"),
  1433 => (x"fa",x"d4",x"ff",x"87"),
  1434 => (x"48",x"66",x"c8",x"87"),
  1435 => (x"c0",x"03",x"a8",x"c7"),
  1436 => (x"e7",x"c2",x"87",x"e5"),
  1437 => (x"78",x"c0",x"48",x"e8"),
  1438 => (x"cb",x"49",x"66",x"c8"),
  1439 => (x"66",x"fc",x"c0",x"91"),
  1440 => (x"4a",x"a1",x"c4",x"81"),
  1441 => (x"52",x"c0",x"4a",x"6a"),
  1442 => (x"48",x"66",x"c8",x"79"),
  1443 => (x"a6",x"cc",x"80",x"c1"),
  1444 => (x"04",x"a8",x"c7",x"58"),
  1445 => (x"ff",x"87",x"db",x"ff"),
  1446 => (x"df",x"ff",x"8e",x"d4"),
  1447 => (x"6f",x"4c",x"87",x"c9"),
  1448 => (x"2a",x"20",x"64",x"61"),
  1449 => (x"3a",x"00",x"20",x"2e"),
  1450 => (x"73",x"1e",x"00",x"20"),
  1451 => (x"9b",x"4b",x"71",x"1e"),
  1452 => (x"c2",x"87",x"c6",x"02"),
  1453 => (x"c0",x"48",x"e4",x"e7"),
  1454 => (x"c2",x"1e",x"c7",x"78"),
  1455 => (x"1e",x"bf",x"e4",x"e7"),
  1456 => (x"1e",x"d9",x"de",x"c1"),
  1457 => (x"bf",x"cc",x"e7",x"c2"),
  1458 => (x"87",x"c1",x"ee",x"49"),
  1459 => (x"e7",x"c2",x"86",x"cc"),
  1460 => (x"e2",x"49",x"bf",x"cc"),
  1461 => (x"9b",x"73",x"87",x"f9"),
  1462 => (x"c1",x"87",x"c8",x"02"),
  1463 => (x"c0",x"49",x"d9",x"de"),
  1464 => (x"ff",x"87",x"c5",x"ef"),
  1465 => (x"1e",x"87",x"c4",x"de"),
  1466 => (x"48",x"c5",x"de",x"c1"),
  1467 => (x"df",x"c1",x"50",x"c0"),
  1468 => (x"ff",x"49",x"bf",x"fc"),
  1469 => (x"c0",x"87",x"c4",x"d9"),
  1470 => (x"1e",x"4f",x"26",x"48"),
  1471 => (x"c1",x"87",x"d3",x"cc"),
  1472 => (x"87",x"e6",x"fe",x"49"),
  1473 => (x"87",x"e8",x"ee",x"fe"),
  1474 => (x"cd",x"02",x"98",x"70"),
  1475 => (x"c2",x"f6",x"fe",x"87"),
  1476 => (x"02",x"98",x"70",x"87"),
  1477 => (x"4a",x"c1",x"87",x"c4"),
  1478 => (x"4a",x"c0",x"87",x"c2"),
  1479 => (x"ce",x"05",x"9a",x"72"),
  1480 => (x"c1",x"1e",x"c0",x"87"),
  1481 => (x"c0",x"49",x"cb",x"dd"),
  1482 => (x"c4",x"87",x"c3",x"fb"),
  1483 => (x"c0",x"87",x"fe",x"86"),
  1484 => (x"d6",x"dd",x"c1",x"1e"),
  1485 => (x"f5",x"fa",x"c0",x"49"),
  1486 => (x"fe",x"1e",x"c0",x"87"),
  1487 => (x"49",x"70",x"87",x"e9"),
  1488 => (x"87",x"ea",x"fa",x"c0"),
  1489 => (x"f8",x"87",x"db",x"c3"),
  1490 => (x"53",x"4f",x"26",x"8e"),
  1491 => (x"61",x"66",x"20",x"44"),
  1492 => (x"64",x"65",x"6c",x"69"),
  1493 => (x"6f",x"42",x"00",x"2e"),
  1494 => (x"6e",x"69",x"74",x"6f"),
  1495 => (x"2e",x"2e",x"2e",x"67"),
  1496 => (x"49",x"c0",x"1e",x"00"),
  1497 => (x"c0",x"87",x"ca",x"d1"),
  1498 => (x"f5",x"87",x"fe",x"f1"),
  1499 => (x"1e",x"4f",x"26",x"87"),
  1500 => (x"48",x"e4",x"e7",x"c2"),
  1501 => (x"e7",x"c2",x"78",x"c0"),
  1502 => (x"78",x"c0",x"48",x"cc"),
  1503 => (x"e0",x"87",x"fc",x"fd"),
  1504 => (x"26",x"48",x"c0",x"87"),
  1505 => (x"01",x"00",x"00",x"4f"),
  1506 => (x"80",x"00",x"00",x"00"),
  1507 => (x"69",x"78",x"45",x"20"),
  1508 => (x"20",x"80",x"00",x"74"),
  1509 => (x"6b",x"63",x"61",x"42"),
  1510 => (x"00",x"0e",x"bd",x"00"),
  1511 => (x"00",x"29",x"f8",x"00"),
  1512 => (x"00",x"00",x"00",x"00"),
  1513 => (x"00",x"00",x"0e",x"bd"),
  1514 => (x"00",x"00",x"2a",x"16"),
  1515 => (x"bd",x"00",x"00",x"00"),
  1516 => (x"34",x"00",x"00",x"0e"),
  1517 => (x"00",x"00",x"00",x"2a"),
  1518 => (x"0e",x"bd",x"00",x"00"),
  1519 => (x"2a",x"52",x"00",x"00"),
  1520 => (x"00",x"00",x"00",x"00"),
  1521 => (x"00",x"0e",x"bd",x"00"),
  1522 => (x"00",x"2a",x"70",x"00"),
  1523 => (x"00",x"00",x"00",x"00"),
  1524 => (x"00",x"00",x"0e",x"bd"),
  1525 => (x"00",x"00",x"2a",x"8e"),
  1526 => (x"bd",x"00",x"00",x"00"),
  1527 => (x"ac",x"00",x"00",x"0e"),
  1528 => (x"00",x"00",x"00",x"2a"),
  1529 => (x"0f",x"70",x"00",x"00"),
  1530 => (x"00",x"00",x"00",x"00"),
  1531 => (x"00",x"00",x"00",x"00"),
  1532 => (x"00",x"11",x"be",x"00"),
  1533 => (x"00",x"00",x"00",x"00"),
  1534 => (x"00",x"00",x"00",x"00"),
  1535 => (x"00",x"00",x"18",x"00"),
  1536 => (x"54",x"4f",x"4f",x"42"),
  1537 => (x"20",x"20",x"20",x"20"),
  1538 => (x"00",x"4d",x"4f",x"52"),
  1539 => (x"48",x"f0",x"fe",x"1e"),
  1540 => (x"09",x"cd",x"78",x"c0"),
  1541 => (x"4f",x"26",x"09",x"79"),
  1542 => (x"f0",x"fe",x"1e",x"1e"),
  1543 => (x"26",x"48",x"7e",x"bf"),
  1544 => (x"fe",x"1e",x"4f",x"26"),
  1545 => (x"78",x"c1",x"48",x"f0"),
  1546 => (x"fe",x"1e",x"4f",x"26"),
  1547 => (x"78",x"c0",x"48",x"f0"),
  1548 => (x"71",x"1e",x"4f",x"26"),
  1549 => (x"7a",x"97",x"c0",x"4a"),
  1550 => (x"c0",x"49",x"a2",x"c1"),
  1551 => (x"49",x"a2",x"ca",x"51"),
  1552 => (x"a2",x"cb",x"51",x"c0"),
  1553 => (x"26",x"51",x"c0",x"49"),
  1554 => (x"5b",x"5e",x"0e",x"4f"),
  1555 => (x"86",x"f0",x"0e",x"5c"),
  1556 => (x"a4",x"ca",x"4c",x"71"),
  1557 => (x"7e",x"69",x"97",x"49"),
  1558 => (x"97",x"4b",x"a4",x"cb"),
  1559 => (x"a6",x"c8",x"48",x"6b"),
  1560 => (x"cc",x"80",x"c1",x"58"),
  1561 => (x"98",x"c7",x"58",x"a6"),
  1562 => (x"6e",x"58",x"a6",x"d0"),
  1563 => (x"a8",x"66",x"cc",x"48"),
  1564 => (x"97",x"87",x"db",x"05"),
  1565 => (x"6b",x"97",x"7e",x"69"),
  1566 => (x"58",x"a6",x"c8",x"48"),
  1567 => (x"a6",x"cc",x"80",x"c1"),
  1568 => (x"d0",x"98",x"c7",x"58"),
  1569 => (x"48",x"6e",x"58",x"a6"),
  1570 => (x"02",x"a8",x"66",x"cc"),
  1571 => (x"d9",x"fe",x"87",x"e5"),
  1572 => (x"4a",x"a4",x"cc",x"87"),
  1573 => (x"72",x"49",x"6b",x"97"),
  1574 => (x"66",x"dc",x"49",x"a1"),
  1575 => (x"7e",x"6b",x"97",x"51"),
  1576 => (x"80",x"c1",x"48",x"6e"),
  1577 => (x"c7",x"58",x"a6",x"c8"),
  1578 => (x"58",x"a6",x"cc",x"98"),
  1579 => (x"c2",x"7b",x"97",x"70"),
  1580 => (x"ed",x"fd",x"87",x"cd"),
  1581 => (x"c2",x"8e",x"f0",x"87"),
  1582 => (x"26",x"4d",x"26",x"87"),
  1583 => (x"26",x"4b",x"26",x"4c"),
  1584 => (x"5b",x"5e",x"0e",x"4f"),
  1585 => (x"f4",x"0e",x"5d",x"5c"),
  1586 => (x"97",x"4d",x"71",x"86"),
  1587 => (x"a5",x"c1",x"7e",x"6d"),
  1588 => (x"48",x"6c",x"97",x"4c"),
  1589 => (x"6e",x"58",x"a6",x"c8"),
  1590 => (x"a8",x"66",x"c4",x"48"),
  1591 => (x"ff",x"87",x"c5",x"05"),
  1592 => (x"87",x"e6",x"c0",x"48"),
  1593 => (x"c2",x"87",x"c3",x"fd"),
  1594 => (x"6c",x"97",x"49",x"a5"),
  1595 => (x"4b",x"a3",x"71",x"4b"),
  1596 => (x"97",x"4b",x"6b",x"97"),
  1597 => (x"48",x"6e",x"7e",x"6c"),
  1598 => (x"a6",x"c8",x"80",x"c1"),
  1599 => (x"cc",x"98",x"c7",x"58"),
  1600 => (x"97",x"70",x"58",x"a6"),
  1601 => (x"87",x"da",x"fc",x"7c"),
  1602 => (x"8e",x"f4",x"48",x"73"),
  1603 => (x"0e",x"87",x"ea",x"fe"),
  1604 => (x"0e",x"5c",x"5b",x"5e"),
  1605 => (x"4c",x"71",x"86",x"f4"),
  1606 => (x"c3",x"4a",x"66",x"d8"),
  1607 => (x"a4",x"c2",x"9a",x"ff"),
  1608 => (x"49",x"6c",x"97",x"4b"),
  1609 => (x"72",x"49",x"a1",x"73"),
  1610 => (x"7e",x"6c",x"97",x"51"),
  1611 => (x"80",x"c1",x"48",x"6e"),
  1612 => (x"c7",x"58",x"a6",x"c8"),
  1613 => (x"58",x"a6",x"cc",x"98"),
  1614 => (x"8e",x"f4",x"54",x"70"),
  1615 => (x"1e",x"87",x"fc",x"fd"),
  1616 => (x"86",x"f4",x"1e",x"73"),
  1617 => (x"e0",x"87",x"e3",x"fb"),
  1618 => (x"c0",x"49",x"4b",x"bf"),
  1619 => (x"02",x"99",x"c0",x"e0"),
  1620 => (x"1e",x"73",x"87",x"cb"),
  1621 => (x"49",x"ca",x"eb",x"c2"),
  1622 => (x"c4",x"87",x"f4",x"fe"),
  1623 => (x"d0",x"49",x"73",x"86"),
  1624 => (x"c1",x"02",x"99",x"c0"),
  1625 => (x"eb",x"c2",x"87",x"c0"),
  1626 => (x"7e",x"bf",x"97",x"d4"),
  1627 => (x"97",x"d5",x"eb",x"c2"),
  1628 => (x"a6",x"c8",x"48",x"bf"),
  1629 => (x"c4",x"48",x"6e",x"58"),
  1630 => (x"c0",x"02",x"a8",x"66"),
  1631 => (x"eb",x"c2",x"87",x"e8"),
  1632 => (x"49",x"bf",x"97",x"d4"),
  1633 => (x"81",x"d6",x"eb",x"c2"),
  1634 => (x"08",x"e0",x"48",x"11"),
  1635 => (x"d4",x"eb",x"c2",x"78"),
  1636 => (x"6e",x"7e",x"bf",x"97"),
  1637 => (x"c8",x"80",x"c1",x"48"),
  1638 => (x"98",x"c7",x"58",x"a6"),
  1639 => (x"c2",x"58",x"a6",x"cc"),
  1640 => (x"c8",x"48",x"d4",x"eb"),
  1641 => (x"bf",x"e4",x"50",x"66"),
  1642 => (x"e0",x"c0",x"49",x"4b"),
  1643 => (x"cb",x"02",x"99",x"c0"),
  1644 => (x"c2",x"1e",x"73",x"87"),
  1645 => (x"fd",x"49",x"de",x"eb"),
  1646 => (x"86",x"c4",x"87",x"d5"),
  1647 => (x"c0",x"d0",x"49",x"73"),
  1648 => (x"c0",x"c1",x"02",x"99"),
  1649 => (x"e8",x"eb",x"c2",x"87"),
  1650 => (x"c2",x"7e",x"bf",x"97"),
  1651 => (x"bf",x"97",x"e9",x"eb"),
  1652 => (x"58",x"a6",x"c8",x"48"),
  1653 => (x"66",x"c4",x"48",x"6e"),
  1654 => (x"e8",x"c0",x"02",x"a8"),
  1655 => (x"e8",x"eb",x"c2",x"87"),
  1656 => (x"c2",x"49",x"bf",x"97"),
  1657 => (x"11",x"81",x"ea",x"eb"),
  1658 => (x"78",x"08",x"e4",x"48"),
  1659 => (x"97",x"e8",x"eb",x"c2"),
  1660 => (x"48",x"6e",x"7e",x"bf"),
  1661 => (x"a6",x"c8",x"80",x"c1"),
  1662 => (x"cc",x"98",x"c7",x"58"),
  1663 => (x"eb",x"c2",x"58",x"a6"),
  1664 => (x"66",x"c8",x"48",x"e8"),
  1665 => (x"87",x"d0",x"f8",x"50"),
  1666 => (x"d5",x"f8",x"7e",x"70"),
  1667 => (x"fa",x"8e",x"f4",x"87"),
  1668 => (x"c2",x"1e",x"87",x"eb"),
  1669 => (x"f8",x"49",x"ca",x"eb"),
  1670 => (x"eb",x"c2",x"87",x"d8"),
  1671 => (x"d1",x"f8",x"49",x"de"),
  1672 => (x"ff",x"e4",x"c1",x"87"),
  1673 => (x"87",x"e4",x"f7",x"49"),
  1674 => (x"26",x"87",x"f7",x"c3"),
  1675 => (x"5b",x"5e",x"0e",x"4f"),
  1676 => (x"71",x"0e",x"5d",x"5c"),
  1677 => (x"ca",x"eb",x"c2",x"4d"),
  1678 => (x"87",x"c5",x"fa",x"49"),
  1679 => (x"b7",x"c0",x"4b",x"70"),
  1680 => (x"c2",x"c3",x"04",x"ab"),
  1681 => (x"ab",x"f0",x"c3",x"87"),
  1682 => (x"c1",x"87",x"c9",x"05"),
  1683 => (x"c1",x"48",x"d1",x"ec"),
  1684 => (x"87",x"e3",x"c2",x"78"),
  1685 => (x"05",x"ab",x"e0",x"c3"),
  1686 => (x"ec",x"c1",x"87",x"c9"),
  1687 => (x"78",x"c1",x"48",x"d5"),
  1688 => (x"c1",x"87",x"d4",x"c2"),
  1689 => (x"02",x"bf",x"d5",x"ec"),
  1690 => (x"c0",x"c2",x"87",x"c6"),
  1691 => (x"87",x"c2",x"4c",x"a3"),
  1692 => (x"ec",x"c1",x"4c",x"73"),
  1693 => (x"c0",x"02",x"bf",x"d1"),
  1694 => (x"49",x"74",x"87",x"e0"),
  1695 => (x"91",x"29",x"b7",x"c4"),
  1696 => (x"81",x"f1",x"ed",x"c1"),
  1697 => (x"9a",x"cf",x"4a",x"74"),
  1698 => (x"48",x"c1",x"92",x"c2"),
  1699 => (x"4a",x"70",x"30",x"72"),
  1700 => (x"48",x"72",x"ba",x"ff"),
  1701 => (x"79",x"70",x"98",x"69"),
  1702 => (x"49",x"74",x"87",x"db"),
  1703 => (x"91",x"29",x"b7",x"c4"),
  1704 => (x"81",x"f1",x"ed",x"c1"),
  1705 => (x"9a",x"cf",x"4a",x"74"),
  1706 => (x"48",x"c3",x"92",x"c2"),
  1707 => (x"4a",x"70",x"30",x"72"),
  1708 => (x"70",x"b0",x"69",x"48"),
  1709 => (x"05",x"9d",x"75",x"79"),
  1710 => (x"ff",x"87",x"f0",x"c0"),
  1711 => (x"e1",x"c8",x"48",x"d0"),
  1712 => (x"48",x"d4",x"ff",x"78"),
  1713 => (x"ec",x"c1",x"78",x"c5"),
  1714 => (x"c3",x"02",x"bf",x"d5"),
  1715 => (x"78",x"e0",x"c3",x"87"),
  1716 => (x"bf",x"d1",x"ec",x"c1"),
  1717 => (x"ff",x"87",x"c6",x"02"),
  1718 => (x"f0",x"c3",x"48",x"d4"),
  1719 => (x"0b",x"d4",x"ff",x"78"),
  1720 => (x"d0",x"ff",x"0b",x"7b"),
  1721 => (x"78",x"e1",x"c8",x"48"),
  1722 => (x"c1",x"78",x"e0",x"c0"),
  1723 => (x"c0",x"48",x"d5",x"ec"),
  1724 => (x"d1",x"ec",x"c1",x"78"),
  1725 => (x"c2",x"78",x"c0",x"48"),
  1726 => (x"f7",x"49",x"ca",x"eb"),
  1727 => (x"4b",x"70",x"87",x"c3"),
  1728 => (x"03",x"ab",x"b7",x"c0"),
  1729 => (x"c0",x"87",x"fe",x"fc"),
  1730 => (x"26",x"4d",x"26",x"48"),
  1731 => (x"26",x"4b",x"26",x"4c"),
  1732 => (x"00",x"00",x"00",x"4f"),
  1733 => (x"00",x"00",x"00",x"00"),
  1734 => (x"4a",x"71",x"1e",x"00"),
  1735 => (x"87",x"cd",x"fc",x"49"),
  1736 => (x"c0",x"1e",x"4f",x"26"),
  1737 => (x"c4",x"49",x"72",x"4a"),
  1738 => (x"f1",x"ed",x"c1",x"91"),
  1739 => (x"c1",x"79",x"c0",x"81"),
  1740 => (x"aa",x"b7",x"d0",x"82"),
  1741 => (x"26",x"87",x"ee",x"04"),
  1742 => (x"5b",x"5e",x"0e",x"4f"),
  1743 => (x"71",x"0e",x"5d",x"5c"),
  1744 => (x"87",x"e6",x"f3",x"4d"),
  1745 => (x"b7",x"c4",x"4a",x"75"),
  1746 => (x"ed",x"c1",x"92",x"2a"),
  1747 => (x"4c",x"75",x"82",x"f1"),
  1748 => (x"94",x"c2",x"9c",x"cf"),
  1749 => (x"74",x"4b",x"49",x"6a"),
  1750 => (x"c2",x"9b",x"c3",x"2b"),
  1751 => (x"70",x"30",x"74",x"48"),
  1752 => (x"74",x"bc",x"ff",x"4c"),
  1753 => (x"70",x"98",x"71",x"48"),
  1754 => (x"87",x"f6",x"f2",x"7a"),
  1755 => (x"d8",x"fe",x"48",x"73"),
  1756 => (x"00",x"00",x"00",x"87"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"5b",x"5e",x"0e",x"00"),
  1773 => (x"4a",x"71",x"0e",x"5c"),
  1774 => (x"87",x"c6",x"02",x"9a"),
  1775 => (x"48",x"ee",x"f5",x"c1"),
  1776 => (x"f5",x"c1",x"78",x"c0"),
  1777 => (x"c0",x"05",x"bf",x"ee"),
  1778 => (x"eb",x"c2",x"87",x"f9"),
  1779 => (x"f0",x"f3",x"49",x"de"),
  1780 => (x"a8",x"b7",x"c0",x"87"),
  1781 => (x"c2",x"87",x"cd",x"04"),
  1782 => (x"f3",x"49",x"de",x"eb"),
  1783 => (x"b7",x"c0",x"87",x"e3"),
  1784 => (x"87",x"f3",x"03",x"a8"),
  1785 => (x"bf",x"ee",x"f5",x"c1"),
  1786 => (x"ee",x"f5",x"c1",x"49"),
  1787 => (x"78",x"a1",x"c1",x"48"),
  1788 => (x"81",x"fe",x"f5",x"c1"),
  1789 => (x"f5",x"c1",x"48",x"11"),
  1790 => (x"f5",x"c1",x"58",x"f6"),
  1791 => (x"78",x"c0",x"48",x"f6"),
  1792 => (x"c1",x"87",x"dc",x"c5"),
  1793 => (x"02",x"bf",x"f6",x"f5"),
  1794 => (x"c2",x"87",x"f2",x"c1"),
  1795 => (x"f2",x"49",x"de",x"eb"),
  1796 => (x"b7",x"c0",x"87",x"ef"),
  1797 => (x"87",x"cd",x"04",x"a8"),
  1798 => (x"bf",x"f6",x"f5",x"c1"),
  1799 => (x"c1",x"88",x"c1",x"48"),
  1800 => (x"db",x"58",x"fa",x"f5"),
  1801 => (x"f2",x"eb",x"c2",x"87"),
  1802 => (x"e8",x"c0",x"49",x"bf"),
  1803 => (x"98",x"70",x"87",x"ed"),
  1804 => (x"c2",x"87",x"cd",x"02"),
  1805 => (x"ef",x"49",x"de",x"eb"),
  1806 => (x"f5",x"c1",x"87",x"f8"),
  1807 => (x"78",x"c0",x"48",x"ee"),
  1808 => (x"bf",x"f2",x"f5",x"c1"),
  1809 => (x"87",x"d7",x"c4",x"05"),
  1810 => (x"bf",x"f6",x"f5",x"c1"),
  1811 => (x"87",x"cf",x"c4",x"05"),
  1812 => (x"bf",x"ee",x"f5",x"c1"),
  1813 => (x"ee",x"f5",x"c1",x"49"),
  1814 => (x"78",x"a1",x"c1",x"48"),
  1815 => (x"81",x"fe",x"f5",x"c1"),
  1816 => (x"c2",x"49",x"4c",x"11"),
  1817 => (x"c0",x"02",x"99",x"c0"),
  1818 => (x"48",x"74",x"87",x"cc"),
  1819 => (x"c1",x"98",x"ff",x"c1"),
  1820 => (x"c3",x"58",x"fa",x"f5"),
  1821 => (x"f5",x"c1",x"87",x"e9"),
  1822 => (x"e2",x"c3",x"5c",x"f6"),
  1823 => (x"f2",x"f5",x"c1",x"87"),
  1824 => (x"fd",x"c0",x"02",x"bf"),
  1825 => (x"ee",x"f5",x"c1",x"87"),
  1826 => (x"f5",x"c1",x"49",x"bf"),
  1827 => (x"a1",x"c1",x"48",x"ee"),
  1828 => (x"fe",x"f5",x"c1",x"78"),
  1829 => (x"49",x"69",x"97",x"81"),
  1830 => (x"de",x"eb",x"c2",x"1e"),
  1831 => (x"87",x"e9",x"ee",x"49"),
  1832 => (x"f5",x"c1",x"86",x"c4"),
  1833 => (x"c1",x"48",x"bf",x"f2"),
  1834 => (x"f6",x"f5",x"c1",x"88"),
  1835 => (x"f6",x"f5",x"c1",x"58"),
  1836 => (x"c0",x"78",x"c1",x"48"),
  1837 => (x"c0",x"49",x"ec",x"f6"),
  1838 => (x"c2",x"87",x"d4",x"e6"),
  1839 => (x"c2",x"58",x"f6",x"eb"),
  1840 => (x"eb",x"c2",x"87",x"dd"),
  1841 => (x"f8",x"ef",x"49",x"de"),
  1842 => (x"c0",x"4b",x"70",x"87"),
  1843 => (x"c2",x"04",x"ab",x"b7"),
  1844 => (x"f5",x"c1",x"87",x"cd"),
  1845 => (x"c0",x"02",x"bf",x"ea"),
  1846 => (x"eb",x"c2",x"87",x"e0"),
  1847 => (x"c0",x"49",x"bf",x"f2"),
  1848 => (x"70",x"87",x"f8",x"e5"),
  1849 => (x"d1",x"c0",x"02",x"98"),
  1850 => (x"c1",x"48",x"c7",x"87"),
  1851 => (x"88",x"bf",x"fa",x"f5"),
  1852 => (x"58",x"fe",x"f5",x"c1"),
  1853 => (x"48",x"ea",x"f5",x"c1"),
  1854 => (x"f5",x"c1",x"78",x"c0"),
  1855 => (x"c1",x"4a",x"bf",x"ea"),
  1856 => (x"f5",x"c1",x"49",x"a2"),
  1857 => (x"eb",x"c2",x"59",x"ee"),
  1858 => (x"52",x"73",x"82",x"f6"),
  1859 => (x"bf",x"fa",x"f5",x"c1"),
  1860 => (x"c0",x"04",x"a9",x"b7"),
  1861 => (x"eb",x"c2",x"87",x"ee"),
  1862 => (x"49",x"bf",x"97",x"f6"),
  1863 => (x"c1",x"49",x"c4",x"1e"),
  1864 => (x"86",x"c4",x"87",x"ec"),
  1865 => (x"97",x"f7",x"eb",x"c2"),
  1866 => (x"d4",x"ff",x"48",x"bf"),
  1867 => (x"eb",x"c2",x"78",x"08"),
  1868 => (x"48",x"bf",x"97",x"f8"),
  1869 => (x"78",x"08",x"d4",x"ff"),
  1870 => (x"c0",x"48",x"d0",x"ff"),
  1871 => (x"f5",x"c1",x"78",x"e0"),
  1872 => (x"78",x"c0",x"48",x"ea"),
  1873 => (x"c0",x"49",x"f4",x"c7"),
  1874 => (x"c2",x"87",x"c4",x"e4"),
  1875 => (x"c2",x"58",x"f6",x"eb"),
  1876 => (x"ed",x"49",x"de",x"eb"),
  1877 => (x"4b",x"70",x"87",x"eb"),
  1878 => (x"03",x"ab",x"b7",x"c0"),
  1879 => (x"c0",x"87",x"f3",x"fd"),
  1880 => (x"4d",x"26",x"87",x"c2"),
  1881 => (x"4b",x"26",x"4c",x"26"),
  1882 => (x"00",x"00",x"4f",x"26"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"00",x"00"),
  1886 => (x"00",x"04",x"00",x"00"),
  1887 => (x"ff",x"01",x"00",x"00"),
  1888 => (x"c8",x"f3",x"08",x"82"),
  1889 => (x"50",x"f3",x"64",x"f3"),
  1890 => (x"01",x"81",x"01",x"f2"),
  1891 => (x"ff",x"1e",x"00",x"f4"),
  1892 => (x"e1",x"c8",x"48",x"d0"),
  1893 => (x"ff",x"48",x"71",x"78"),
  1894 => (x"c4",x"78",x"08",x"d4"),
  1895 => (x"d4",x"ff",x"48",x"66"),
  1896 => (x"4f",x"26",x"78",x"08"),
  1897 => (x"c4",x"4a",x"71",x"1e"),
  1898 => (x"72",x"1e",x"49",x"66"),
  1899 => (x"87",x"de",x"ff",x"49"),
  1900 => (x"c0",x"48",x"d0",x"ff"),
  1901 => (x"26",x"26",x"78",x"e0"),
  1902 => (x"1e",x"73",x"1e",x"4f"),
  1903 => (x"66",x"c8",x"4b",x"71"),
  1904 => (x"4a",x"73",x"1e",x"49"),
  1905 => (x"49",x"a2",x"e0",x"c1"),
  1906 => (x"26",x"87",x"d9",x"ff"),
  1907 => (x"4d",x"26",x"87",x"c4"),
  1908 => (x"4b",x"26",x"4c",x"26"),
  1909 => (x"ff",x"1e",x"4f",x"26"),
  1910 => (x"ff",x"c3",x"4a",x"d4"),
  1911 => (x"48",x"d0",x"ff",x"7a"),
  1912 => (x"de",x"78",x"e1",x"c0"),
  1913 => (x"fa",x"eb",x"c2",x"7a"),
  1914 => (x"48",x"49",x"7a",x"bf"),
  1915 => (x"7a",x"70",x"28",x"c8"),
  1916 => (x"28",x"d0",x"48",x"71"),
  1917 => (x"48",x"71",x"7a",x"70"),
  1918 => (x"7a",x"70",x"28",x"d8"),
  1919 => (x"c0",x"48",x"d0",x"ff"),
  1920 => (x"4f",x"26",x"78",x"e0"),
  1921 => (x"48",x"d0",x"ff",x"1e"),
  1922 => (x"71",x"78",x"c9",x"c8"),
  1923 => (x"08",x"d4",x"ff",x"48"),
  1924 => (x"1e",x"4f",x"26",x"78"),
  1925 => (x"eb",x"49",x"4a",x"71"),
  1926 => (x"48",x"d0",x"ff",x"87"),
  1927 => (x"4f",x"26",x"78",x"c8"),
  1928 => (x"71",x"1e",x"73",x"1e"),
  1929 => (x"ca",x"ec",x"c2",x"4b"),
  1930 => (x"87",x"c3",x"02",x"bf"),
  1931 => (x"ff",x"87",x"eb",x"c2"),
  1932 => (x"c9",x"c8",x"48",x"d0"),
  1933 => (x"c0",x"48",x"73",x"78"),
  1934 => (x"d4",x"ff",x"b0",x"e0"),
  1935 => (x"eb",x"c2",x"78",x"08"),
  1936 => (x"78",x"c0",x"48",x"fe"),
  1937 => (x"c5",x"02",x"66",x"c8"),
  1938 => (x"49",x"ff",x"c3",x"87"),
  1939 => (x"49",x"c0",x"87",x"c2"),
  1940 => (x"59",x"c6",x"ec",x"c2"),
  1941 => (x"c6",x"02",x"66",x"cc"),
  1942 => (x"d5",x"d5",x"c5",x"87"),
  1943 => (x"cf",x"87",x"c4",x"4a"),
  1944 => (x"c2",x"4a",x"ff",x"ff"),
  1945 => (x"c2",x"5a",x"ca",x"ec"),
  1946 => (x"c1",x"48",x"ca",x"ec"),
  1947 => (x"26",x"87",x"c4",x"78"),
  1948 => (x"26",x"4c",x"26",x"4d"),
  1949 => (x"0e",x"4f",x"26",x"4b"),
  1950 => (x"5d",x"5c",x"5b",x"5e"),
  1951 => (x"c2",x"4a",x"71",x"0e"),
  1952 => (x"4c",x"bf",x"c6",x"ec"),
  1953 => (x"cb",x"02",x"9a",x"72"),
  1954 => (x"91",x"c8",x"49",x"87"),
  1955 => (x"4b",x"d6",x"f8",x"c1"),
  1956 => (x"87",x"c4",x"83",x"71"),
  1957 => (x"4b",x"d6",x"fc",x"c1"),
  1958 => (x"49",x"13",x"4d",x"c0"),
  1959 => (x"ec",x"c2",x"99",x"74"),
  1960 => (x"71",x"48",x"bf",x"c2"),
  1961 => (x"08",x"d4",x"ff",x"b8"),
  1962 => (x"2c",x"b7",x"c1",x"78"),
  1963 => (x"ad",x"b7",x"c8",x"85"),
  1964 => (x"c2",x"87",x"e7",x"04"),
  1965 => (x"48",x"bf",x"fe",x"eb"),
  1966 => (x"ec",x"c2",x"80",x"c8"),
  1967 => (x"ee",x"fe",x"58",x"c2"),
  1968 => (x"1e",x"73",x"1e",x"87"),
  1969 => (x"4a",x"13",x"4b",x"71"),
  1970 => (x"87",x"cb",x"02",x"9a"),
  1971 => (x"e6",x"fe",x"49",x"72"),
  1972 => (x"9a",x"4a",x"13",x"87"),
  1973 => (x"fe",x"87",x"f5",x"05"),
  1974 => (x"c2",x"1e",x"87",x"d9"),
  1975 => (x"49",x"bf",x"fe",x"eb"),
  1976 => (x"48",x"fe",x"eb",x"c2"),
  1977 => (x"c4",x"78",x"a1",x"c1"),
  1978 => (x"03",x"a9",x"b7",x"c0"),
  1979 => (x"d4",x"ff",x"87",x"db"),
  1980 => (x"c2",x"ec",x"c2",x"48"),
  1981 => (x"eb",x"c2",x"78",x"bf"),
  1982 => (x"c2",x"49",x"bf",x"fe"),
  1983 => (x"c1",x"48",x"fe",x"eb"),
  1984 => (x"c0",x"c4",x"78",x"a1"),
  1985 => (x"e5",x"04",x"a9",x"b7"),
  1986 => (x"48",x"d0",x"ff",x"87"),
  1987 => (x"ec",x"c2",x"78",x"c8"),
  1988 => (x"78",x"c0",x"48",x"ca"),
  1989 => (x"00",x"00",x"4f",x"26"),
  1990 => (x"00",x"00",x"00",x"00"),
  1991 => (x"00",x"00",x"00",x"00"),
  1992 => (x"00",x"5f",x"5f",x"00"),
  1993 => (x"03",x"00",x"00",x"00"),
  1994 => (x"03",x"03",x"00",x"03"),
  1995 => (x"7f",x"14",x"00",x"00"),
  1996 => (x"7f",x"7f",x"14",x"7f"),
  1997 => (x"24",x"00",x"00",x"14"),
  1998 => (x"3a",x"6b",x"6b",x"2e"),
  1999 => (x"6a",x"4c",x"00",x"12"),
  2000 => (x"56",x"6c",x"18",x"36"),
  2001 => (x"7e",x"30",x"00",x"32"),
  2002 => (x"3a",x"77",x"59",x"4f"),
  2003 => (x"00",x"00",x"40",x"68"),
  2004 => (x"00",x"03",x"07",x"04"),
  2005 => (x"00",x"00",x"00",x"00"),
  2006 => (x"41",x"63",x"3e",x"1c"),
  2007 => (x"00",x"00",x"00",x"00"),
  2008 => (x"1c",x"3e",x"63",x"41"),
  2009 => (x"2a",x"08",x"00",x"00"),
  2010 => (x"3e",x"1c",x"1c",x"3e"),
  2011 => (x"08",x"00",x"08",x"2a"),
  2012 => (x"08",x"3e",x"3e",x"08"),
  2013 => (x"00",x"00",x"00",x"08"),
  2014 => (x"00",x"60",x"e0",x"80"),
  2015 => (x"08",x"00",x"00",x"00"),
  2016 => (x"08",x"08",x"08",x"08"),
  2017 => (x"00",x"00",x"00",x"08"),
  2018 => (x"00",x"60",x"60",x"00"),
  2019 => (x"60",x"40",x"00",x"00"),
  2020 => (x"06",x"0c",x"18",x"30"),
  2021 => (x"3e",x"00",x"01",x"03"),
  2022 => (x"7f",x"4d",x"59",x"7f"),
  2023 => (x"04",x"00",x"00",x"3e"),
  2024 => (x"00",x"7f",x"7f",x"06"),
  2025 => (x"42",x"00",x"00",x"00"),
  2026 => (x"4f",x"59",x"71",x"63"),
  2027 => (x"22",x"00",x"00",x"46"),
  2028 => (x"7f",x"49",x"49",x"63"),
  2029 => (x"1c",x"18",x"00",x"36"),
  2030 => (x"7f",x"7f",x"13",x"16"),
  2031 => (x"27",x"00",x"00",x"10"),
  2032 => (x"7d",x"45",x"45",x"67"),
  2033 => (x"3c",x"00",x"00",x"39"),
  2034 => (x"79",x"49",x"4b",x"7e"),
  2035 => (x"01",x"00",x"00",x"30"),
  2036 => (x"0f",x"79",x"71",x"01"),
  2037 => (x"36",x"00",x"00",x"07"),
  2038 => (x"7f",x"49",x"49",x"7f"),
  2039 => (x"06",x"00",x"00",x"36"),
  2040 => (x"3f",x"69",x"49",x"4f"),
  2041 => (x"00",x"00",x"00",x"1e"),
  2042 => (x"00",x"66",x"66",x"00"),
  2043 => (x"00",x"00",x"00",x"00"),
  2044 => (x"00",x"66",x"e6",x"80"),
  2045 => (x"08",x"00",x"00",x"00"),
  2046 => (x"22",x"14",x"14",x"08"),
  2047 => (x"14",x"00",x"00",x"22"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

