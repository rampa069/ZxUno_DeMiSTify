library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e4ecc287",
    12 => x"86c0c84e",
    13 => x"49e4ecc2",
    14 => x"48f4d9c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e4dc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c348724c",
    72 => x"7c7098ff",
    73 => x"bff4d9c2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"29d04966",
    81 => x"ffc34871",
    82 => x"d07c7098",
    83 => x"29c84966",
    84 => x"ffc34871",
    85 => x"d07c7098",
    86 => x"ffc34866",
    87 => x"727c7098",
    88 => x"7129d049",
    89 => x"98ffc348",
    90 => x"4b6c7c70",
    91 => x"4dfff0c9",
    92 => x"05abffc3",
    93 => x"ffc387d0",
    94 => x"c14b6c7c",
    95 => x"87c6028d",
    96 => x"02abffc3",
    97 => x"487387f0",
    98 => x"1e87fffd",
    99 => x"d4ff49c0",
   100 => x"78ffc348",
   101 => x"c8c381c1",
   102 => x"f104a9b7",
   103 => x"1e4f2687",
   104 => x"87e71e73",
   105 => x"4bdff8c4",
   106 => x"ffc01ec0",
   107 => x"49f7c1f0",
   108 => x"c487dffd",
   109 => x"05a8c186",
   110 => x"ff87eac0",
   111 => x"ffc348d4",
   112 => x"c0c0c178",
   113 => x"1ec0c0c0",
   114 => x"c1f0e1c0",
   115 => x"c1fd49e9",
   116 => x"7086c487",
   117 => x"87ca0598",
   118 => x"c348d4ff",
   119 => x"48c178ff",
   120 => x"e6fe87cb",
   121 => x"058bc187",
   122 => x"c087fdfe",
   123 => x"87defc48",
   124 => x"ff1e731e",
   125 => x"ffc348d4",
   126 => x"c04bd378",
   127 => x"f0ffc01e",
   128 => x"fc49c1c1",
   129 => x"86c487cc",
   130 => x"ca059870",
   131 => x"48d4ff87",
   132 => x"c178ffc3",
   133 => x"fd87cb48",
   134 => x"8bc187f1",
   135 => x"87dbff05",
   136 => x"e9fb48c0",
   137 => x"5b5e0e87",
   138 => x"d4ff0e5c",
   139 => x"87dbfd4c",
   140 => x"c01eeac6",
   141 => x"c8c1f0e1",
   142 => x"87d6fb49",
   143 => x"a8c186c4",
   144 => x"fe87c802",
   145 => x"48c087ea",
   146 => x"fa87e2c1",
   147 => x"497087d2",
   148 => x"99ffffcf",
   149 => x"02a9eac6",
   150 => x"d3fe87c8",
   151 => x"c148c087",
   152 => x"ffc387cb",
   153 => x"4bf1c07c",
   154 => x"7087f4fc",
   155 => x"ebc00298",
   156 => x"c01ec087",
   157 => x"fac1f0ff",
   158 => x"87d6fa49",
   159 => x"987086c4",
   160 => x"c387d905",
   161 => x"496c7cff",
   162 => x"7c7cffc3",
   163 => x"c0c17c7c",
   164 => x"87c40299",
   165 => x"87d548c1",
   166 => x"87d148c0",
   167 => x"c405abc2",
   168 => x"c848c087",
   169 => x"058bc187",
   170 => x"c087fdfe",
   171 => x"87dcf948",
   172 => x"c21e731e",
   173 => x"c148f4d9",
   174 => x"ff4bc778",
   175 => x"78c248d0",
   176 => x"ff87c8fb",
   177 => x"78c348d0",
   178 => x"e5c01ec0",
   179 => x"49c0c1d0",
   180 => x"c487fff8",
   181 => x"05a8c186",
   182 => x"c24b87c1",
   183 => x"87c505ab",
   184 => x"f9c048c0",
   185 => x"058bc187",
   186 => x"fc87d0ff",
   187 => x"d9c287f7",
   188 => x"987058f8",
   189 => x"c187cd05",
   190 => x"f0ffc01e",
   191 => x"f849d0c1",
   192 => x"86c487d0",
   193 => x"c348d4ff",
   194 => x"fdc278ff",
   195 => x"fcd9c287",
   196 => x"48d0ff58",
   197 => x"d4ff78c2",
   198 => x"78ffc348",
   199 => x"edf748c1",
   200 => x"5b5e0e87",
   201 => x"710e5d5c",
   202 => x"c54cc04b",
   203 => x"4adfcdee",
   204 => x"c348d4ff",
   205 => x"486878ff",
   206 => x"05a8fec3",
   207 => x"ff87fec0",
   208 => x"9b734dd4",
   209 => x"d087cc02",
   210 => x"49731e66",
   211 => x"c487e8f5",
   212 => x"ff87d686",
   213 => x"d1c448d0",
   214 => x"7dffc378",
   215 => x"c14866d0",
   216 => x"58a6d488",
   217 => x"f0059870",
   218 => x"48d4ff87",
   219 => x"7878ffc3",
   220 => x"c5059b73",
   221 => x"48d0ff87",
   222 => x"4ac178d0",
   223 => x"058ac14c",
   224 => x"7487edfe",
   225 => x"87c2f648",
   226 => x"711e731e",
   227 => x"ff4bc04a",
   228 => x"ffc348d4",
   229 => x"48d0ff78",
   230 => x"ff78c3c4",
   231 => x"ffc348d4",
   232 => x"c01e7278",
   233 => x"d1c1f0ff",
   234 => x"87e6f549",
   235 => x"987086c4",
   236 => x"c887d205",
   237 => x"66cc1ec0",
   238 => x"87e5fd49",
   239 => x"4b7086c4",
   240 => x"c248d0ff",
   241 => x"f5487378",
   242 => x"5e0e87c4",
   243 => x"0e5d5c5b",
   244 => x"ffc01ec0",
   245 => x"49c9c1f0",
   246 => x"d287f7f4",
   247 => x"fcd9c21e",
   248 => x"87fdfc49",
   249 => x"4cc086c8",
   250 => x"b7d284c1",
   251 => x"87f804ac",
   252 => x"97fcd9c2",
   253 => x"c0c349bf",
   254 => x"a9c0c199",
   255 => x"87e7c005",
   256 => x"97c3dac2",
   257 => x"31d049bf",
   258 => x"97c4dac2",
   259 => x"32c84abf",
   260 => x"dac2b172",
   261 => x"4abf97c5",
   262 => x"cf4c71b1",
   263 => x"9cffffff",
   264 => x"34ca84c1",
   265 => x"c287e7c1",
   266 => x"bf97c5da",
   267 => x"c631c149",
   268 => x"c6dac299",
   269 => x"c74abf97",
   270 => x"b1722ab7",
   271 => x"97c1dac2",
   272 => x"cf4d4abf",
   273 => x"c2dac29d",
   274 => x"c34abf97",
   275 => x"c232ca9a",
   276 => x"bf97c3da",
   277 => x"7333c24b",
   278 => x"c4dac2b2",
   279 => x"c34bbf97",
   280 => x"b7c69bc0",
   281 => x"c2b2732b",
   282 => x"7148c181",
   283 => x"c1497030",
   284 => x"70307548",
   285 => x"c14c724d",
   286 => x"c8947184",
   287 => x"06adb7c0",
   288 => x"34c187cc",
   289 => x"c0c82db7",
   290 => x"ff01adb7",
   291 => x"487487f4",
   292 => x"0e87f7f1",
   293 => x"5d5c5b5e",
   294 => x"c286f80e",
   295 => x"c048e2e2",
   296 => x"dadac278",
   297 => x"fb49c01e",
   298 => x"86c487de",
   299 => x"c5059870",
   300 => x"c948c087",
   301 => x"4dc087c0",
   302 => x"edc07ec1",
   303 => x"c249bfe6",
   304 => x"714ad0db",
   305 => x"e0ee4bc8",
   306 => x"05987087",
   307 => x"7ec087c2",
   308 => x"bfe2edc0",
   309 => x"ecdbc249",
   310 => x"4bc8714a",
   311 => x"7087caee",
   312 => x"87c20598",
   313 => x"026e7ec0",
   314 => x"c287fdc0",
   315 => x"4dbfe0e1",
   316 => x"9fd8e2c2",
   317 => x"c5487ebf",
   318 => x"05a8ead6",
   319 => x"e1c287c7",
   320 => x"ce4dbfe0",
   321 => x"ca486e87",
   322 => x"02a8d5e9",
   323 => x"48c087c5",
   324 => x"c287e3c7",
   325 => x"751edada",
   326 => x"87ecf949",
   327 => x"987086c4",
   328 => x"c087c505",
   329 => x"87cec748",
   330 => x"bfe2edc0",
   331 => x"ecdbc249",
   332 => x"4bc8714a",
   333 => x"7087f2ec",
   334 => x"87c80598",
   335 => x"48e2e2c2",
   336 => x"87da78c1",
   337 => x"bfe6edc0",
   338 => x"d0dbc249",
   339 => x"4bc8714a",
   340 => x"7087d6ec",
   341 => x"c5c00298",
   342 => x"c648c087",
   343 => x"e2c287d8",
   344 => x"49bf97d8",
   345 => x"05a9d5c1",
   346 => x"c287cdc0",
   347 => x"bf97d9e2",
   348 => x"a9eac249",
   349 => x"87c5c002",
   350 => x"f9c548c0",
   351 => x"dadac287",
   352 => x"487ebf97",
   353 => x"02a8e9c3",
   354 => x"6e87cec0",
   355 => x"a8ebc348",
   356 => x"87c5c002",
   357 => x"ddc548c0",
   358 => x"e5dac287",
   359 => x"9949bf97",
   360 => x"87ccc005",
   361 => x"97e6dac2",
   362 => x"a9c249bf",
   363 => x"87c5c002",
   364 => x"c1c548c0",
   365 => x"e7dac287",
   366 => x"c248bf97",
   367 => x"7058dee2",
   368 => x"88c1484c",
   369 => x"58e2e2c2",
   370 => x"97e8dac2",
   371 => x"817549bf",
   372 => x"97e9dac2",
   373 => x"32c84abf",
   374 => x"c27ea172",
   375 => x"6e48efe6",
   376 => x"eadac278",
   377 => x"c848bf97",
   378 => x"e2c258a6",
   379 => x"c202bfe2",
   380 => x"edc087cf",
   381 => x"c249bfe2",
   382 => x"714aecdb",
   383 => x"e8e94bc8",
   384 => x"02987087",
   385 => x"c087c5c0",
   386 => x"87eac348",
   387 => x"bfdae2c2",
   388 => x"c3e7c24c",
   389 => x"ffdac25c",
   390 => x"c849bf97",
   391 => x"fedac231",
   392 => x"a14abf97",
   393 => x"c0dbc249",
   394 => x"d04abf97",
   395 => x"49a17232",
   396 => x"97c1dbc2",
   397 => x"32d84abf",
   398 => x"c449a172",
   399 => x"e6c29166",
   400 => x"c281bfef",
   401 => x"c259f7e6",
   402 => x"bf97c7db",
   403 => x"c232c84a",
   404 => x"bf97c6db",
   405 => x"c24aa24b",
   406 => x"bf97c8db",
   407 => x"7333d04b",
   408 => x"dbc24aa2",
   409 => x"4bbf97c9",
   410 => x"33d89bcf",
   411 => x"c24aa273",
   412 => x"c25afbe6",
   413 => x"c292748a",
   414 => x"7248fbe6",
   415 => x"c1c178a1",
   416 => x"ecdac287",
   417 => x"c849bf97",
   418 => x"ebdac231",
   419 => x"a14abf97",
   420 => x"c731c549",
   421 => x"29c981ff",
   422 => x"59c3e7c2",
   423 => x"97f1dac2",
   424 => x"32c84abf",
   425 => x"97f0dac2",
   426 => x"4aa24bbf",
   427 => x"6e9266c4",
   428 => x"ffe6c282",
   429 => x"f7e6c25a",
   430 => x"c278c048",
   431 => x"7248f3e6",
   432 => x"e7c278a1",
   433 => x"e6c248c3",
   434 => x"c278bff7",
   435 => x"c248c7e7",
   436 => x"78bffbe6",
   437 => x"bfe2e2c2",
   438 => x"87c9c002",
   439 => x"30c44874",
   440 => x"c9c07e70",
   441 => x"ffe6c287",
   442 => x"30c448bf",
   443 => x"e2c27e70",
   444 => x"786e48e6",
   445 => x"8ef848c1",
   446 => x"4c264d26",
   447 => x"4f264b26",
   448 => x"5c5b5e0e",
   449 => x"4a710e5d",
   450 => x"bfe2e2c2",
   451 => x"7287cb02",
   452 => x"722bc74b",
   453 => x"9dffc14d",
   454 => x"4b7287c9",
   455 => x"4d722bc8",
   456 => x"c29dffc3",
   457 => x"83bfefe6",
   458 => x"bfdeedc0",
   459 => x"87d902ab",
   460 => x"5be2edc0",
   461 => x"1edadac2",
   462 => x"cbf14973",
   463 => x"7086c487",
   464 => x"87c50598",
   465 => x"e6c048c0",
   466 => x"e2e2c287",
   467 => x"87d202bf",
   468 => x"91c44975",
   469 => x"81dadac2",
   470 => x"ffcf4c69",
   471 => x"9cffffff",
   472 => x"497587cb",
   473 => x"dac291c2",
   474 => x"699f81da",
   475 => x"fe48744c",
   476 => x"5e0e87c6",
   477 => x"0e5d5c5b",
   478 => x"4c7186f8",
   479 => x"87c5059c",
   480 => x"c0c348c0",
   481 => x"7ea4c887",
   482 => x"d878c048",
   483 => x"87c70266",
   484 => x"bf9766d8",
   485 => x"c087c505",
   486 => x"87e9c248",
   487 => x"49c11ec0",
   488 => x"87e3c749",
   489 => x"4d7086c4",
   490 => x"c2c1029d",
   491 => x"eae2c287",
   492 => x"4966d84a",
   493 => x"7087d7e2",
   494 => x"f2c00298",
   495 => x"d84a7587",
   496 => x"4bcb4966",
   497 => x"7087fce2",
   498 => x"e2c00298",
   499 => x"751ec087",
   500 => x"87c7029d",
   501 => x"c048a6c8",
   502 => x"c887c578",
   503 => x"78c148a6",
   504 => x"c64966c8",
   505 => x"86c487e1",
   506 => x"059d4d70",
   507 => x"7587fefe",
   508 => x"cec1029d",
   509 => x"49a5dc87",
   510 => x"7869486e",
   511 => x"c449a5da",
   512 => x"a4c448a6",
   513 => x"48699f78",
   514 => x"780866c4",
   515 => x"bfe2e2c2",
   516 => x"d487d202",
   517 => x"699f49a5",
   518 => x"ffffc049",
   519 => x"d0487199",
   520 => x"c27e7030",
   521 => x"6e7ec087",
   522 => x"bf66c448",
   523 => x"0866c480",
   524 => x"cc7cc078",
   525 => x"66c449a4",
   526 => x"a4d079bf",
   527 => x"c179c049",
   528 => x"c087c248",
   529 => x"fa8ef848",
   530 => x"5e0e87ee",
   531 => x"710e5c5b",
   532 => x"c1029c4c",
   533 => x"a4c887cb",
   534 => x"c1026949",
   535 => x"496c87c3",
   536 => x"714866cc",
   537 => x"58a6d080",
   538 => x"e2c2b970",
   539 => x"ff4abfde",
   540 => x"719972ba",
   541 => x"e5c00299",
   542 => x"4ba4c487",
   543 => x"fff9496b",
   544 => x"c27b7087",
   545 => x"49bfdae2",
   546 => x"7c71816c",
   547 => x"c2b966cc",
   548 => x"4abfdee2",
   549 => x"9972baff",
   550 => x"ff059971",
   551 => x"66cc87db",
   552 => x"87d6f97c",
   553 => x"711e731e",
   554 => x"c7029b4b",
   555 => x"49a3c887",
   556 => x"87c50569",
   557 => x"f6c048c0",
   558 => x"f3e6c287",
   559 => x"a3c449bf",
   560 => x"c24a6a4a",
   561 => x"dae2c28a",
   562 => x"a17292bf",
   563 => x"dee2c249",
   564 => x"9a6b4abf",
   565 => x"c049a172",
   566 => x"c859e2ed",
   567 => x"ea711e66",
   568 => x"86c487e6",
   569 => x"c4059870",
   570 => x"c248c087",
   571 => x"f848c187",
   572 => x"731e87ca",
   573 => x"9b4b711e",
   574 => x"87e4c002",
   575 => x"5bc7e7c2",
   576 => x"8ac24a73",
   577 => x"bfdae2c2",
   578 => x"e6c29249",
   579 => x"7248bff3",
   580 => x"cbe7c280",
   581 => x"c4487158",
   582 => x"eae2c230",
   583 => x"87edc058",
   584 => x"48c3e7c2",
   585 => x"bff7e6c2",
   586 => x"c7e7c278",
   587 => x"fbe6c248",
   588 => x"e2c278bf",
   589 => x"c902bfe2",
   590 => x"dae2c287",
   591 => x"31c449bf",
   592 => x"e6c287c7",
   593 => x"c449bfff",
   594 => x"eae2c231",
   595 => x"87ecf659",
   596 => x"5c5b5e0e",
   597 => x"c04a710e",
   598 => x"029a724b",
   599 => x"da87e0c0",
   600 => x"699f49a2",
   601 => x"e2e2c24b",
   602 => x"87cf02bf",
   603 => x"9f49a2d4",
   604 => x"c04c4969",
   605 => x"d09cffff",
   606 => x"c087c234",
   607 => x"73b3744c",
   608 => x"87eefd49",
   609 => x"0e87f3f5",
   610 => x"5d5c5b5e",
   611 => x"7186f40e",
   612 => x"727ec04a",
   613 => x"87d8029a",
   614 => x"48d6dac2",
   615 => x"dac278c0",
   616 => x"e7c248ce",
   617 => x"c278bfc7",
   618 => x"c248d2da",
   619 => x"78bfc3e7",
   620 => x"48f7e2c2",
   621 => x"e2c250c0",
   622 => x"c249bfe6",
   623 => x"4abfd6da",
   624 => x"c403aa71",
   625 => x"497287c9",
   626 => x"c00599cf",
   627 => x"edc087e9",
   628 => x"dac248de",
   629 => x"c278bfce",
   630 => x"c21edada",
   631 => x"49bfceda",
   632 => x"48cedac2",
   633 => x"7178a1c1",
   634 => x"c487dde6",
   635 => x"daedc086",
   636 => x"dadac248",
   637 => x"c087cc78",
   638 => x"48bfdaed",
   639 => x"c080e0c0",
   640 => x"c258deed",
   641 => x"48bfd6da",
   642 => x"dac280c1",
   643 => x"5a2758da",
   644 => x"bf00000b",
   645 => x"9d4dbf97",
   646 => x"87e3c202",
   647 => x"02ade5c3",
   648 => x"c087dcc2",
   649 => x"4bbfdaed",
   650 => x"1149a3cb",
   651 => x"05accf4c",
   652 => x"7587d2c1",
   653 => x"c199df49",
   654 => x"c291cd89",
   655 => x"c181eae2",
   656 => x"51124aa3",
   657 => x"124aa3c3",
   658 => x"4aa3c551",
   659 => x"a3c75112",
   660 => x"c951124a",
   661 => x"51124aa3",
   662 => x"124aa3ce",
   663 => x"4aa3d051",
   664 => x"a3d25112",
   665 => x"d451124a",
   666 => x"51124aa3",
   667 => x"124aa3d6",
   668 => x"4aa3d851",
   669 => x"a3dc5112",
   670 => x"de51124a",
   671 => x"51124aa3",
   672 => x"fac07ec1",
   673 => x"c8497487",
   674 => x"ebc00599",
   675 => x"d0497487",
   676 => x"87d10599",
   677 => x"c00266dc",
   678 => x"497387cb",
   679 => x"700f66dc",
   680 => x"d3c00298",
   681 => x"c0056e87",
   682 => x"e2c287c6",
   683 => x"50c048ea",
   684 => x"bfdaedc0",
   685 => x"87ddc248",
   686 => x"48f7e2c2",
   687 => x"c27e50c0",
   688 => x"49bfe6e2",
   689 => x"bfd6dac2",
   690 => x"04aa714a",
   691 => x"c287f7fb",
   692 => x"05bfc7e7",
   693 => x"c287c8c0",
   694 => x"02bfe2e2",
   695 => x"c287f4c1",
   696 => x"49bfd2da",
   697 => x"c287d9f0",
   698 => x"c458d6da",
   699 => x"dac248a6",
   700 => x"c278bfd2",
   701 => x"02bfe2e2",
   702 => x"c487d8c0",
   703 => x"ffcf4966",
   704 => x"99f8ffff",
   705 => x"c5c002a9",
   706 => x"c04cc087",
   707 => x"4cc187e1",
   708 => x"c487dcc0",
   709 => x"ffcf4966",
   710 => x"02a999f8",
   711 => x"c887c8c0",
   712 => x"78c048a6",
   713 => x"c887c5c0",
   714 => x"78c148a6",
   715 => x"744c66c8",
   716 => x"dec0059c",
   717 => x"4966c487",
   718 => x"e2c289c2",
   719 => x"c291bfda",
   720 => x"48bff3e6",
   721 => x"dac28071",
   722 => x"dac258d2",
   723 => x"78c048d6",
   724 => x"c087e3f9",
   725 => x"ee8ef448",
   726 => x"000087de",
   727 => x"ffff0000",
   728 => x"0b6affff",
   729 => x"0b730000",
   730 => x"41460000",
   731 => x"20323354",
   732 => x"46002020",
   733 => x"36315441",
   734 => x"00202020",
   735 => x"48d4ff1e",
   736 => x"6878ffc3",
   737 => x"1e4f2648",
   738 => x"c348d4ff",
   739 => x"d0ff78ff",
   740 => x"78e1c048",
   741 => x"d448d4ff",
   742 => x"cbe7c278",
   743 => x"bfd4ff48",
   744 => x"1e4f2650",
   745 => x"c048d0ff",
   746 => x"4f2678e0",
   747 => x"87ccff1e",
   748 => x"02994970",
   749 => x"fbc087c6",
   750 => x"87f105a9",
   751 => x"4f264871",
   752 => x"5c5b5e0e",
   753 => x"c04b710e",
   754 => x"87f0fe4c",
   755 => x"02994970",
   756 => x"c087f9c0",
   757 => x"c002a9ec",
   758 => x"fbc087f2",
   759 => x"ebc002a9",
   760 => x"b766cc87",
   761 => x"87c703ac",
   762 => x"c20266d0",
   763 => x"71537187",
   764 => x"87c20299",
   765 => x"c3fe84c1",
   766 => x"99497087",
   767 => x"c087cd02",
   768 => x"c702a9ec",
   769 => x"a9fbc087",
   770 => x"87d5ff05",
   771 => x"c30266d0",
   772 => x"7b97c087",
   773 => x"05a9ecc0",
   774 => x"4a7487c4",
   775 => x"4a7487c5",
   776 => x"728a0ac0",
   777 => x"2687c248",
   778 => x"264c264d",
   779 => x"1e4f264b",
   780 => x"7087c9fd",
   781 => x"aaf0c04a",
   782 => x"c087c904",
   783 => x"c301aaf9",
   784 => x"8af0c087",
   785 => x"04aac1c1",
   786 => x"dac187c9",
   787 => x"87c301aa",
   788 => x"728af7c0",
   789 => x"0e4f2648",
   790 => x"0e5c5b5e",
   791 => x"d4ff4a71",
   792 => x"c049724b",
   793 => x"4c7087e7",
   794 => x"87c2029c",
   795 => x"d0ff8cc1",
   796 => x"c178c548",
   797 => x"49747bd5",
   798 => x"dec131c6",
   799 => x"4abf97c5",
   800 => x"70b07148",
   801 => x"48d0ff7b",
   802 => x"dcfe78c4",
   803 => x"5b5e0e87",
   804 => x"f80e5d5c",
   805 => x"c04c7186",
   806 => x"87ebfb7e",
   807 => x"f4c04bc0",
   808 => x"49bf97fa",
   809 => x"cf04a9c0",
   810 => x"87c0fc87",
   811 => x"f4c083c1",
   812 => x"49bf97fa",
   813 => x"87f106ab",
   814 => x"97faf4c0",
   815 => x"87cf02bf",
   816 => x"7087f9fa",
   817 => x"c6029949",
   818 => x"a9ecc087",
   819 => x"c087f105",
   820 => x"87e8fa4b",
   821 => x"e3fa4d70",
   822 => x"58a6c887",
   823 => x"7087ddfa",
   824 => x"c883c14a",
   825 => x"699749a4",
   826 => x"c702ad49",
   827 => x"adffc087",
   828 => x"87e7c005",
   829 => x"9749a4c9",
   830 => x"66c44969",
   831 => x"87c702a9",
   832 => x"a8ffc048",
   833 => x"ca87d405",
   834 => x"699749a4",
   835 => x"c602aa49",
   836 => x"aaffc087",
   837 => x"c187c405",
   838 => x"c087d07e",
   839 => x"c602adec",
   840 => x"adfbc087",
   841 => x"c087c405",
   842 => x"6e7ec14b",
   843 => x"87e1fe02",
   844 => x"7387f0f9",
   845 => x"fb8ef848",
   846 => x"0e0087ed",
   847 => x"5d5c5b5e",
   848 => x"7186f80e",
   849 => x"4bd4ff4d",
   850 => x"e7c21e75",
   851 => x"e1e849d0",
   852 => x"7086c487",
   853 => x"cac40298",
   854 => x"48a6c487",
   855 => x"bfc7dec1",
   856 => x"fb497578",
   857 => x"d0ff87f1",
   858 => x"c178c548",
   859 => x"4ac07bd6",
   860 => x"1149a275",
   861 => x"cb82c17b",
   862 => x"f304aab7",
   863 => x"c34acc87",
   864 => x"82c17bff",
   865 => x"aab7e0c0",
   866 => x"ff87f404",
   867 => x"78c448d0",
   868 => x"c57bffc3",
   869 => x"7bd3c178",
   870 => x"78c47bc1",
   871 => x"b7c04866",
   872 => x"eec206a8",
   873 => x"d8e7c287",
   874 => x"66c44cbf",
   875 => x"c8887448",
   876 => x"9c7458a6",
   877 => x"87f7c102",
   878 => x"7edadac2",
   879 => x"8c4dc0c8",
   880 => x"03acb7c0",
   881 => x"c0c887c6",
   882 => x"4cc04da4",
   883 => x"97cbe7c2",
   884 => x"99d049bf",
   885 => x"c087d002",
   886 => x"d0e7c21e",
   887 => x"87c4eb49",
   888 => x"4a7086c4",
   889 => x"c287edc0",
   890 => x"c21edada",
   891 => x"ea49d0e7",
   892 => x"86c487f2",
   893 => x"d0ff4a70",
   894 => x"78c5c848",
   895 => x"6e7bd4c1",
   896 => x"6e7bbf97",
   897 => x"7080c148",
   898 => x"058dc17e",
   899 => x"ff87f0ff",
   900 => x"78c448d0",
   901 => x"c5059a72",
   902 => x"c148c087",
   903 => x"1ec187c7",
   904 => x"49d0e7c2",
   905 => x"c487e3e8",
   906 => x"059c7486",
   907 => x"c487c9fe",
   908 => x"b7c04866",
   909 => x"87d106a8",
   910 => x"48d0e7c2",
   911 => x"80d078c0",
   912 => x"80f478c0",
   913 => x"bfdce7c2",
   914 => x"4866c478",
   915 => x"01a8b7c0",
   916 => x"ff87d2fd",
   917 => x"78c548d0",
   918 => x"c07bd3c1",
   919 => x"c178c47b",
   920 => x"c087c248",
   921 => x"268ef848",
   922 => x"264c264d",
   923 => x"0e4f264b",
   924 => x"5d5c5b5e",
   925 => x"4b711e0e",
   926 => x"ab4d4cc0",
   927 => x"87e8c004",
   928 => x"1ecdf2c0",
   929 => x"c4029d75",
   930 => x"c24ac087",
   931 => x"724ac187",
   932 => x"87f3eb49",
   933 => x"7e7086c4",
   934 => x"056e84c1",
   935 => x"4c7387c2",
   936 => x"ac7385c1",
   937 => x"87d8ff06",
   938 => x"fe26486e",
   939 => x"711e87f9",
   940 => x"0566c44a",
   941 => x"497287c5",
   942 => x"2687c0fa",
   943 => x"5b5e0e4f",
   944 => x"1e0e5d5c",
   945 => x"de494c71",
   946 => x"f8e7c291",
   947 => x"9785714d",
   948 => x"dcc1026d",
   949 => x"e4e7c287",
   950 => x"817449bf",
   951 => x"87cffe71",
   952 => x"98487e70",
   953 => x"87f2c002",
   954 => x"4bece7c2",
   955 => x"49cb4a70",
   956 => x"87f3c6ff",
   957 => x"93cb4b74",
   958 => x"83d9dec1",
   959 => x"fcc083c4",
   960 => x"49747bf5",
   961 => x"87cecdc1",
   962 => x"dec17b75",
   963 => x"49bf97c6",
   964 => x"ece7c21e",
   965 => x"87d6fe49",
   966 => x"497486c4",
   967 => x"87f6ccc1",
   968 => x"cec149c0",
   969 => x"e7c287d5",
   970 => x"78c048cc",
   971 => x"f9dd49c1",
   972 => x"f2fc2687",
   973 => x"616f4c87",
   974 => x"676e6964",
   975 => x"002e2e2e",
   976 => x"711e731e",
   977 => x"e7c2494a",
   978 => x"7181bfe4",
   979 => x"7087e0fc",
   980 => x"c4029b4b",
   981 => x"f7e74987",
   982 => x"e4e7c287",
   983 => x"c178c048",
   984 => x"87c6dd49",
   985 => x"1e87c4fc",
   986 => x"cdc149c0",
   987 => x"4f2687cd",
   988 => x"494a711e",
   989 => x"dec191cb",
   990 => x"81c881d9",
   991 => x"e7c24811",
   992 => x"e7c258d0",
   993 => x"78c048e4",
   994 => x"dddc49c1",
   995 => x"1e4f2687",
   996 => x"d2029971",
   997 => x"eedfc187",
   998 => x"f750c048",
   999 => x"f0fdc080",
  1000 => x"d2dec140",
  1001 => x"c187ce78",
  1002 => x"c148eadf",
  1003 => x"fc78cbde",
  1004 => x"e7fdc080",
  1005 => x"0e4f2678",
  1006 => x"5d5c5b5e",
  1007 => x"c286f40e",
  1008 => x"c04ddada",
  1009 => x"48a6c44c",
  1010 => x"e7c278c0",
  1011 => x"c048bfe4",
  1012 => x"c0c106a8",
  1013 => x"dadac287",
  1014 => x"c0029848",
  1015 => x"f2c087f7",
  1016 => x"66c81ecd",
  1017 => x"c487c702",
  1018 => x"78c048a6",
  1019 => x"a6c487c5",
  1020 => x"c478c148",
  1021 => x"cee64966",
  1022 => x"7086c487",
  1023 => x"c484c14d",
  1024 => x"80c14866",
  1025 => x"c258a6c8",
  1026 => x"acbfe4e7",
  1027 => x"7587c603",
  1028 => x"c9ff059d",
  1029 => x"754cc087",
  1030 => x"dcc3029d",
  1031 => x"cdf2c087",
  1032 => x"0266c81e",
  1033 => x"a6cc87c7",
  1034 => x"c578c048",
  1035 => x"48a6cc87",
  1036 => x"66cc78c1",
  1037 => x"87cfe549",
  1038 => x"7e7086c4",
  1039 => x"c2029848",
  1040 => x"cb4987e4",
  1041 => x"49699781",
  1042 => x"c10299d0",
  1043 => x"497487d4",
  1044 => x"dec191cb",
  1045 => x"fdc081d9",
  1046 => x"81c879c0",
  1047 => x"7451ffc3",
  1048 => x"c291de49",
  1049 => x"714df8e7",
  1050 => x"97c1c285",
  1051 => x"49a5c17d",
  1052 => x"c251e0c0",
  1053 => x"bf97eae2",
  1054 => x"c187d202",
  1055 => x"4ba5c284",
  1056 => x"4aeae2c2",
  1057 => x"c0ff49db",
  1058 => x"d9c187dd",
  1059 => x"49a5cd87",
  1060 => x"84c151c0",
  1061 => x"6e4ba5c2",
  1062 => x"ff49cb4a",
  1063 => x"c187c8c0",
  1064 => x"497487c4",
  1065 => x"dec191cb",
  1066 => x"fac081d9",
  1067 => x"e2c279fd",
  1068 => x"02bf97ea",
  1069 => x"497487d8",
  1070 => x"84c191de",
  1071 => x"4bf8e7c2",
  1072 => x"e2c28371",
  1073 => x"49dd4aea",
  1074 => x"87dbfffe",
  1075 => x"4b7487d8",
  1076 => x"e7c293de",
  1077 => x"a3cb83f8",
  1078 => x"c151c049",
  1079 => x"4a6e7384",
  1080 => x"fffe49cb",
  1081 => x"66c487c1",
  1082 => x"c880c148",
  1083 => x"acc758a6",
  1084 => x"87c5c003",
  1085 => x"e4fc056e",
  1086 => x"f4487487",
  1087 => x"87e7f58e",
  1088 => x"711e731e",
  1089 => x"91cb494b",
  1090 => x"81d9dec1",
  1091 => x"c14aa1c8",
  1092 => x"1248c5de",
  1093 => x"4aa1c950",
  1094 => x"48faf4c0",
  1095 => x"81ca5012",
  1096 => x"48c6dec1",
  1097 => x"dec15011",
  1098 => x"49bf97c6",
  1099 => x"f549c01e",
  1100 => x"e7c287fc",
  1101 => x"78de48cc",
  1102 => x"edd549c1",
  1103 => x"eaf42687",
  1104 => x"5b5e0e87",
  1105 => x"f40e5d5c",
  1106 => x"494d7186",
  1107 => x"dec191cb",
  1108 => x"a1c881d9",
  1109 => x"7ea1ca4a",
  1110 => x"c248a6c4",
  1111 => x"78bffaeb",
  1112 => x"4bbf976e",
  1113 => x"734c66c4",
  1114 => x"cc48122c",
  1115 => x"9c7058a6",
  1116 => x"81c984c1",
  1117 => x"b7496997",
  1118 => x"87c204ac",
  1119 => x"976e4cc0",
  1120 => x"66c84abf",
  1121 => x"ff317249",
  1122 => x"9966c4b9",
  1123 => x"30724874",
  1124 => x"71484a70",
  1125 => x"feebc2b0",
  1126 => x"f9f0c058",
  1127 => x"d449c087",
  1128 => x"497587c8",
  1129 => x"87eec2c1",
  1130 => x"faf28ef4",
  1131 => x"1e731e87",
  1132 => x"fe494b71",
  1133 => x"497387cb",
  1134 => x"f287c6fe",
  1135 => x"731e87ed",
  1136 => x"c64b711e",
  1137 => x"db024aa3",
  1138 => x"028ac187",
  1139 => x"028a87d6",
  1140 => x"8a87dac1",
  1141 => x"87fcc002",
  1142 => x"e1c0028a",
  1143 => x"cb028a87",
  1144 => x"87dbc187",
  1145 => x"c7f649c7",
  1146 => x"87dec187",
  1147 => x"bfe4e7c2",
  1148 => x"87cbc102",
  1149 => x"c288c148",
  1150 => x"c158e8e7",
  1151 => x"e7c287c1",
  1152 => x"c002bfe8",
  1153 => x"e7c287f9",
  1154 => x"c148bfe4",
  1155 => x"e8e7c280",
  1156 => x"87ebc058",
  1157 => x"bfe4e7c2",
  1158 => x"c289c649",
  1159 => x"c059e8e7",
  1160 => x"da03a9b7",
  1161 => x"e4e7c287",
  1162 => x"d278c048",
  1163 => x"e8e7c287",
  1164 => x"87cb02bf",
  1165 => x"bfe4e7c2",
  1166 => x"c280c648",
  1167 => x"c058e8e7",
  1168 => x"87e6d149",
  1169 => x"c0c14973",
  1170 => x"def087cc",
  1171 => x"5b5e0e87",
  1172 => x"ff0e5d5c",
  1173 => x"a6dc86d4",
  1174 => x"48a6c859",
  1175 => x"80c478c0",
  1176 => x"7866c0c1",
  1177 => x"78c180c4",
  1178 => x"78c180c4",
  1179 => x"48e8e7c2",
  1180 => x"e7c278c1",
  1181 => x"de48bfcc",
  1182 => x"87c905a8",
  1183 => x"cc87f8f4",
  1184 => x"e4cf58a6",
  1185 => x"87ffe387",
  1186 => x"e387e1e4",
  1187 => x"4c7087ee",
  1188 => x"02acfbc0",
  1189 => x"d887fbc1",
  1190 => x"edc10566",
  1191 => x"66fcc087",
  1192 => x"6a82c44a",
  1193 => x"c11e727e",
  1194 => x"c448deda",
  1195 => x"a1c84966",
  1196 => x"7141204a",
  1197 => x"87f905aa",
  1198 => x"4a265110",
  1199 => x"4866fcc0",
  1200 => x"78c0c4c1",
  1201 => x"81c7496a",
  1202 => x"fcc05174",
  1203 => x"81c84966",
  1204 => x"fcc051c1",
  1205 => x"81c94966",
  1206 => x"fcc051c0",
  1207 => x"81ca4966",
  1208 => x"1ec151c0",
  1209 => x"496a1ed8",
  1210 => x"d3e381c8",
  1211 => x"c186c887",
  1212 => x"c04866c0",
  1213 => x"87c701a8",
  1214 => x"c148a6c8",
  1215 => x"c187ce78",
  1216 => x"c14866c0",
  1217 => x"58a6d088",
  1218 => x"dfe287c3",
  1219 => x"48a6d087",
  1220 => x"9c7478c2",
  1221 => x"87cdcd02",
  1222 => x"c14866c8",
  1223 => x"03a866c4",
  1224 => x"dc87c2cd",
  1225 => x"78c048a6",
  1226 => x"78c080e8",
  1227 => x"7087cde1",
  1228 => x"acd0c14c",
  1229 => x"87d5c205",
  1230 => x"e37e66c4",
  1231 => x"a6c887f1",
  1232 => x"87f8e058",
  1233 => x"ecc04c70",
  1234 => x"ebc105ac",
  1235 => x"4966c887",
  1236 => x"fcc091cb",
  1237 => x"a1c48166",
  1238 => x"c84d6a4a",
  1239 => x"66c44aa1",
  1240 => x"f0fdc052",
  1241 => x"87d4e079",
  1242 => x"029c4c70",
  1243 => x"fbc087d8",
  1244 => x"87d202ac",
  1245 => x"c3e05574",
  1246 => x"9c4c7087",
  1247 => x"c087c702",
  1248 => x"ff05acfb",
  1249 => x"e0c087ee",
  1250 => x"55c1c255",
  1251 => x"d87d97c0",
  1252 => x"a86e4866",
  1253 => x"c887db05",
  1254 => x"66cc4866",
  1255 => x"87ca04a8",
  1256 => x"c14866c8",
  1257 => x"58a6cc80",
  1258 => x"66cc87c8",
  1259 => x"d088c148",
  1260 => x"dfff58a6",
  1261 => x"4c7087c6",
  1262 => x"05acd0c1",
  1263 => x"66d487c8",
  1264 => x"d880c148",
  1265 => x"d0c158a6",
  1266 => x"ebfd02ac",
  1267 => x"4866c487",
  1268 => x"05a866d8",
  1269 => x"c087e0c9",
  1270 => x"c048a6e0",
  1271 => x"c0487478",
  1272 => x"7e7088fb",
  1273 => x"c9029848",
  1274 => x"cb4887e2",
  1275 => x"487e7088",
  1276 => x"cdc10298",
  1277 => x"88c94887",
  1278 => x"98487e70",
  1279 => x"87fec302",
  1280 => x"7088c448",
  1281 => x"0298487e",
  1282 => x"c14887ce",
  1283 => x"487e7088",
  1284 => x"e9c30298",
  1285 => x"87d6c887",
  1286 => x"c048a6dc",
  1287 => x"ddff78f0",
  1288 => x"4c7087da",
  1289 => x"02acecc0",
  1290 => x"c087c4c0",
  1291 => x"c05ca6e0",
  1292 => x"cd02acec",
  1293 => x"c3ddff87",
  1294 => x"c04c7087",
  1295 => x"ff05acec",
  1296 => x"ecc087f3",
  1297 => x"c4c002ac",
  1298 => x"efdcff87",
  1299 => x"ca1ec087",
  1300 => x"4966d01e",
  1301 => x"c4c191cb",
  1302 => x"80714866",
  1303 => x"c858a6cc",
  1304 => x"80c44866",
  1305 => x"cc58a6d0",
  1306 => x"ff49bf66",
  1307 => x"c187d1dd",
  1308 => x"d41ede1e",
  1309 => x"ff49bf66",
  1310 => x"d087c5dd",
  1311 => x"48497086",
  1312 => x"c08808c0",
  1313 => x"c058a6e8",
  1314 => x"eec006a8",
  1315 => x"66e4c087",
  1316 => x"03a8dd48",
  1317 => x"c487e4c0",
  1318 => x"c049bf66",
  1319 => x"c08166e4",
  1320 => x"e4c051e0",
  1321 => x"81c14966",
  1322 => x"81bf66c4",
  1323 => x"c051c1c2",
  1324 => x"c24966e4",
  1325 => x"bf66c481",
  1326 => x"6e51c081",
  1327 => x"c0c4c148",
  1328 => x"c8496e78",
  1329 => x"5166d081",
  1330 => x"81c9496e",
  1331 => x"6e5166d4",
  1332 => x"dc81ca49",
  1333 => x"66d05166",
  1334 => x"d480c148",
  1335 => x"66c858a6",
  1336 => x"a866cc48",
  1337 => x"87cbc004",
  1338 => x"c14866c8",
  1339 => x"58a6cc80",
  1340 => x"cc87d9c5",
  1341 => x"88c14866",
  1342 => x"c558a6d0",
  1343 => x"dcff87ce",
  1344 => x"e8c087ed",
  1345 => x"dcff58a6",
  1346 => x"e0c087e5",
  1347 => x"ecc058a6",
  1348 => x"cac005a8",
  1349 => x"48a6dc87",
  1350 => x"7866e4c0",
  1351 => x"ff87c4c0",
  1352 => x"c887d9d9",
  1353 => x"91cb4966",
  1354 => x"4866fcc0",
  1355 => x"7e708071",
  1356 => x"6e82c84a",
  1357 => x"c081ca49",
  1358 => x"dc5166e4",
  1359 => x"81c14966",
  1360 => x"8966e4c0",
  1361 => x"307148c1",
  1362 => x"89c14970",
  1363 => x"c27a9771",
  1364 => x"49bffaeb",
  1365 => x"2966e4c0",
  1366 => x"484a6a97",
  1367 => x"ecc09871",
  1368 => x"496e58a6",
  1369 => x"4d6981c4",
  1370 => x"c44866d8",
  1371 => x"c002a866",
  1372 => x"a6c487c8",
  1373 => x"c078c048",
  1374 => x"a6c487c5",
  1375 => x"c478c148",
  1376 => x"e0c01e66",
  1377 => x"ff49751e",
  1378 => x"c887f5d8",
  1379 => x"c04c7086",
  1380 => x"c106acb7",
  1381 => x"857487d4",
  1382 => x"7449e0c0",
  1383 => x"c14b7589",
  1384 => x"714ae7da",
  1385 => x"87ffebfe",
  1386 => x"e0c085c2",
  1387 => x"80c14866",
  1388 => x"58a6e4c0",
  1389 => x"4966e8c0",
  1390 => x"a97081c1",
  1391 => x"87c8c002",
  1392 => x"c048a6c4",
  1393 => x"87c5c078",
  1394 => x"c148a6c4",
  1395 => x"1e66c478",
  1396 => x"c049a4c2",
  1397 => x"887148e0",
  1398 => x"751e4970",
  1399 => x"dfd7ff49",
  1400 => x"c086c887",
  1401 => x"ff01a8b7",
  1402 => x"e0c087c0",
  1403 => x"d1c00266",
  1404 => x"c9496e87",
  1405 => x"66e0c081",
  1406 => x"c1486e51",
  1407 => x"c078c1c5",
  1408 => x"496e87cc",
  1409 => x"51c281c9",
  1410 => x"c6c1486e",
  1411 => x"66c878ed",
  1412 => x"a866cc48",
  1413 => x"87cbc004",
  1414 => x"c14866c8",
  1415 => x"58a6cc80",
  1416 => x"cc87e9c0",
  1417 => x"88c14866",
  1418 => x"c058a6d0",
  1419 => x"d5ff87de",
  1420 => x"4c7087fa",
  1421 => x"c187d5c0",
  1422 => x"c005acc6",
  1423 => x"66d087c8",
  1424 => x"d480c148",
  1425 => x"d5ff58a6",
  1426 => x"4c7087e2",
  1427 => x"c14866d4",
  1428 => x"58a6d880",
  1429 => x"c0029c74",
  1430 => x"66c887cb",
  1431 => x"66c4c148",
  1432 => x"fef204a8",
  1433 => x"fad4ff87",
  1434 => x"4866c887",
  1435 => x"c003a8c7",
  1436 => x"e7c287e5",
  1437 => x"78c048e8",
  1438 => x"cb4966c8",
  1439 => x"66fcc091",
  1440 => x"4aa1c481",
  1441 => x"52c04a6a",
  1442 => x"4866c879",
  1443 => x"a6cc80c1",
  1444 => x"04a8c758",
  1445 => x"ff87dbff",
  1446 => x"dfff8ed4",
  1447 => x"6f4c87c9",
  1448 => x"2a206461",
  1449 => x"3a00202e",
  1450 => x"731e0020",
  1451 => x"9b4b711e",
  1452 => x"c287c602",
  1453 => x"c048e4e7",
  1454 => x"c21ec778",
  1455 => x"1ebfe4e7",
  1456 => x"1ed9dec1",
  1457 => x"bfcce7c2",
  1458 => x"87c1ee49",
  1459 => x"e7c286cc",
  1460 => x"e249bfcc",
  1461 => x"9b7387f9",
  1462 => x"c187c802",
  1463 => x"c049d9de",
  1464 => x"ff87c5ef",
  1465 => x"1e87c4de",
  1466 => x"48c5dec1",
  1467 => x"dfc150c0",
  1468 => x"ff49bffc",
  1469 => x"c087c4d9",
  1470 => x"1e4f2648",
  1471 => x"c187d3cc",
  1472 => x"87e6fe49",
  1473 => x"87e8eefe",
  1474 => x"cd029870",
  1475 => x"c2f6fe87",
  1476 => x"02987087",
  1477 => x"4ac187c4",
  1478 => x"4ac087c2",
  1479 => x"ce059a72",
  1480 => x"c11ec087",
  1481 => x"c049cbdd",
  1482 => x"c487c3fb",
  1483 => x"c087fe86",
  1484 => x"d6ddc11e",
  1485 => x"f5fac049",
  1486 => x"fe1ec087",
  1487 => x"497087e9",
  1488 => x"87eafac0",
  1489 => x"f887dbc3",
  1490 => x"534f268e",
  1491 => x"61662044",
  1492 => x"64656c69",
  1493 => x"6f42002e",
  1494 => x"6e69746f",
  1495 => x"2e2e2e67",
  1496 => x"49c01e00",
  1497 => x"c087cad1",
  1498 => x"f587fef1",
  1499 => x"1e4f2687",
  1500 => x"48e4e7c2",
  1501 => x"e7c278c0",
  1502 => x"78c048cc",
  1503 => x"e087fcfd",
  1504 => x"2648c087",
  1505 => x"0100004f",
  1506 => x"80000000",
  1507 => x"69784520",
  1508 => x"20800074",
  1509 => x"6b636142",
  1510 => x"000ebd00",
  1511 => x"0029f800",
  1512 => x"00000000",
  1513 => x"00000ebd",
  1514 => x"00002a16",
  1515 => x"bd000000",
  1516 => x"3400000e",
  1517 => x"0000002a",
  1518 => x"0ebd0000",
  1519 => x"2a520000",
  1520 => x"00000000",
  1521 => x"000ebd00",
  1522 => x"002a7000",
  1523 => x"00000000",
  1524 => x"00000ebd",
  1525 => x"00002a8e",
  1526 => x"bd000000",
  1527 => x"ac00000e",
  1528 => x"0000002a",
  1529 => x"0f700000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"0011be00",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00001800",
  1536 => x"544f4f42",
  1537 => x"20202020",
  1538 => x"004d4f52",
  1539 => x"48f0fe1e",
  1540 => x"09cd78c0",
  1541 => x"4f260979",
  1542 => x"f0fe1e1e",
  1543 => x"26487ebf",
  1544 => x"fe1e4f26",
  1545 => x"78c148f0",
  1546 => x"fe1e4f26",
  1547 => x"78c048f0",
  1548 => x"711e4f26",
  1549 => x"7a97c04a",
  1550 => x"c049a2c1",
  1551 => x"49a2ca51",
  1552 => x"a2cb51c0",
  1553 => x"2651c049",
  1554 => x"5b5e0e4f",
  1555 => x"86f00e5c",
  1556 => x"a4ca4c71",
  1557 => x"7e699749",
  1558 => x"974ba4cb",
  1559 => x"a6c8486b",
  1560 => x"cc80c158",
  1561 => x"98c758a6",
  1562 => x"6e58a6d0",
  1563 => x"a866cc48",
  1564 => x"9787db05",
  1565 => x"6b977e69",
  1566 => x"58a6c848",
  1567 => x"a6cc80c1",
  1568 => x"d098c758",
  1569 => x"486e58a6",
  1570 => x"02a866cc",
  1571 => x"d9fe87e5",
  1572 => x"4aa4cc87",
  1573 => x"72496b97",
  1574 => x"66dc49a1",
  1575 => x"7e6b9751",
  1576 => x"80c1486e",
  1577 => x"c758a6c8",
  1578 => x"58a6cc98",
  1579 => x"c27b9770",
  1580 => x"edfd87cd",
  1581 => x"c28ef087",
  1582 => x"264d2687",
  1583 => x"264b264c",
  1584 => x"5b5e0e4f",
  1585 => x"f40e5d5c",
  1586 => x"974d7186",
  1587 => x"a5c17e6d",
  1588 => x"486c974c",
  1589 => x"6e58a6c8",
  1590 => x"a866c448",
  1591 => x"ff87c505",
  1592 => x"87e6c048",
  1593 => x"c287c3fd",
  1594 => x"6c9749a5",
  1595 => x"4ba3714b",
  1596 => x"974b6b97",
  1597 => x"486e7e6c",
  1598 => x"a6c880c1",
  1599 => x"cc98c758",
  1600 => x"977058a6",
  1601 => x"87dafc7c",
  1602 => x"8ef44873",
  1603 => x"0e87eafe",
  1604 => x"0e5c5b5e",
  1605 => x"4c7186f4",
  1606 => x"c34a66d8",
  1607 => x"a4c29aff",
  1608 => x"496c974b",
  1609 => x"7249a173",
  1610 => x"7e6c9751",
  1611 => x"80c1486e",
  1612 => x"c758a6c8",
  1613 => x"58a6cc98",
  1614 => x"8ef45470",
  1615 => x"1e87fcfd",
  1616 => x"86f41e73",
  1617 => x"e087e3fb",
  1618 => x"c0494bbf",
  1619 => x"0299c0e0",
  1620 => x"1e7387cb",
  1621 => x"49caebc2",
  1622 => x"c487f4fe",
  1623 => x"d0497386",
  1624 => x"c10299c0",
  1625 => x"ebc287c0",
  1626 => x"7ebf97d4",
  1627 => x"97d5ebc2",
  1628 => x"a6c848bf",
  1629 => x"c4486e58",
  1630 => x"c002a866",
  1631 => x"ebc287e8",
  1632 => x"49bf97d4",
  1633 => x"81d6ebc2",
  1634 => x"08e04811",
  1635 => x"d4ebc278",
  1636 => x"6e7ebf97",
  1637 => x"c880c148",
  1638 => x"98c758a6",
  1639 => x"c258a6cc",
  1640 => x"c848d4eb",
  1641 => x"bfe45066",
  1642 => x"e0c0494b",
  1643 => x"cb0299c0",
  1644 => x"c21e7387",
  1645 => x"fd49deeb",
  1646 => x"86c487d5",
  1647 => x"c0d04973",
  1648 => x"c0c10299",
  1649 => x"e8ebc287",
  1650 => x"c27ebf97",
  1651 => x"bf97e9eb",
  1652 => x"58a6c848",
  1653 => x"66c4486e",
  1654 => x"e8c002a8",
  1655 => x"e8ebc287",
  1656 => x"c249bf97",
  1657 => x"1181eaeb",
  1658 => x"7808e448",
  1659 => x"97e8ebc2",
  1660 => x"486e7ebf",
  1661 => x"a6c880c1",
  1662 => x"cc98c758",
  1663 => x"ebc258a6",
  1664 => x"66c848e8",
  1665 => x"87d0f850",
  1666 => x"d5f87e70",
  1667 => x"fa8ef487",
  1668 => x"c21e87eb",
  1669 => x"f849caeb",
  1670 => x"ebc287d8",
  1671 => x"d1f849de",
  1672 => x"ffe4c187",
  1673 => x"87e4f749",
  1674 => x"2687f7c3",
  1675 => x"5b5e0e4f",
  1676 => x"710e5d5c",
  1677 => x"caebc24d",
  1678 => x"87c5fa49",
  1679 => x"b7c04b70",
  1680 => x"c2c304ab",
  1681 => x"abf0c387",
  1682 => x"c187c905",
  1683 => x"c148d1ec",
  1684 => x"87e3c278",
  1685 => x"05abe0c3",
  1686 => x"ecc187c9",
  1687 => x"78c148d5",
  1688 => x"c187d4c2",
  1689 => x"02bfd5ec",
  1690 => x"c0c287c6",
  1691 => x"87c24ca3",
  1692 => x"ecc14c73",
  1693 => x"c002bfd1",
  1694 => x"497487e0",
  1695 => x"9129b7c4",
  1696 => x"81f1edc1",
  1697 => x"9acf4a74",
  1698 => x"48c192c2",
  1699 => x"4a703072",
  1700 => x"4872baff",
  1701 => x"79709869",
  1702 => x"497487db",
  1703 => x"9129b7c4",
  1704 => x"81f1edc1",
  1705 => x"9acf4a74",
  1706 => x"48c392c2",
  1707 => x"4a703072",
  1708 => x"70b06948",
  1709 => x"059d7579",
  1710 => x"ff87f0c0",
  1711 => x"e1c848d0",
  1712 => x"48d4ff78",
  1713 => x"ecc178c5",
  1714 => x"c302bfd5",
  1715 => x"78e0c387",
  1716 => x"bfd1ecc1",
  1717 => x"ff87c602",
  1718 => x"f0c348d4",
  1719 => x"0bd4ff78",
  1720 => x"d0ff0b7b",
  1721 => x"78e1c848",
  1722 => x"c178e0c0",
  1723 => x"c048d5ec",
  1724 => x"d1ecc178",
  1725 => x"c278c048",
  1726 => x"f749caeb",
  1727 => x"4b7087c3",
  1728 => x"03abb7c0",
  1729 => x"c087fefc",
  1730 => x"264d2648",
  1731 => x"264b264c",
  1732 => x"0000004f",
  1733 => x"00000000",
  1734 => x"4a711e00",
  1735 => x"87cdfc49",
  1736 => x"c01e4f26",
  1737 => x"c449724a",
  1738 => x"f1edc191",
  1739 => x"c179c081",
  1740 => x"aab7d082",
  1741 => x"2687ee04",
  1742 => x"5b5e0e4f",
  1743 => x"710e5d5c",
  1744 => x"87e6f34d",
  1745 => x"b7c44a75",
  1746 => x"edc1922a",
  1747 => x"4c7582f1",
  1748 => x"94c29ccf",
  1749 => x"744b496a",
  1750 => x"c29bc32b",
  1751 => x"70307448",
  1752 => x"74bcff4c",
  1753 => x"70987148",
  1754 => x"87f6f27a",
  1755 => x"d8fe4873",
  1756 => x"00000087",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"5b5e0e00",
  1773 => x"4a710e5c",
  1774 => x"87c6029a",
  1775 => x"48eef5c1",
  1776 => x"f5c178c0",
  1777 => x"c005bfee",
  1778 => x"ebc287f9",
  1779 => x"f0f349de",
  1780 => x"a8b7c087",
  1781 => x"c287cd04",
  1782 => x"f349deeb",
  1783 => x"b7c087e3",
  1784 => x"87f303a8",
  1785 => x"bfeef5c1",
  1786 => x"eef5c149",
  1787 => x"78a1c148",
  1788 => x"81fef5c1",
  1789 => x"f5c14811",
  1790 => x"f5c158f6",
  1791 => x"78c048f6",
  1792 => x"c187dcc5",
  1793 => x"02bff6f5",
  1794 => x"c287f2c1",
  1795 => x"f249deeb",
  1796 => x"b7c087ef",
  1797 => x"87cd04a8",
  1798 => x"bff6f5c1",
  1799 => x"c188c148",
  1800 => x"db58faf5",
  1801 => x"f2ebc287",
  1802 => x"e8c049bf",
  1803 => x"987087ed",
  1804 => x"c287cd02",
  1805 => x"ef49deeb",
  1806 => x"f5c187f8",
  1807 => x"78c048ee",
  1808 => x"bff2f5c1",
  1809 => x"87d7c405",
  1810 => x"bff6f5c1",
  1811 => x"87cfc405",
  1812 => x"bfeef5c1",
  1813 => x"eef5c149",
  1814 => x"78a1c148",
  1815 => x"81fef5c1",
  1816 => x"c2494c11",
  1817 => x"c00299c0",
  1818 => x"487487cc",
  1819 => x"c198ffc1",
  1820 => x"c358faf5",
  1821 => x"f5c187e9",
  1822 => x"e2c35cf6",
  1823 => x"f2f5c187",
  1824 => x"fdc002bf",
  1825 => x"eef5c187",
  1826 => x"f5c149bf",
  1827 => x"a1c148ee",
  1828 => x"fef5c178",
  1829 => x"49699781",
  1830 => x"deebc21e",
  1831 => x"87e9ee49",
  1832 => x"f5c186c4",
  1833 => x"c148bff2",
  1834 => x"f6f5c188",
  1835 => x"f6f5c158",
  1836 => x"c078c148",
  1837 => x"c049ecf6",
  1838 => x"c287d4e6",
  1839 => x"c258f6eb",
  1840 => x"ebc287dd",
  1841 => x"f8ef49de",
  1842 => x"c04b7087",
  1843 => x"c204abb7",
  1844 => x"f5c187cd",
  1845 => x"c002bfea",
  1846 => x"ebc287e0",
  1847 => x"c049bff2",
  1848 => x"7087f8e5",
  1849 => x"d1c00298",
  1850 => x"c148c787",
  1851 => x"88bffaf5",
  1852 => x"58fef5c1",
  1853 => x"48eaf5c1",
  1854 => x"f5c178c0",
  1855 => x"c14abfea",
  1856 => x"f5c149a2",
  1857 => x"ebc259ee",
  1858 => x"527382f6",
  1859 => x"bffaf5c1",
  1860 => x"c004a9b7",
  1861 => x"ebc287ee",
  1862 => x"49bf97f6",
  1863 => x"c149c41e",
  1864 => x"86c487ec",
  1865 => x"97f7ebc2",
  1866 => x"d4ff48bf",
  1867 => x"ebc27808",
  1868 => x"48bf97f8",
  1869 => x"7808d4ff",
  1870 => x"c048d0ff",
  1871 => x"f5c178e0",
  1872 => x"78c048ea",
  1873 => x"c049f4c7",
  1874 => x"c287c4e4",
  1875 => x"c258f6eb",
  1876 => x"ed49deeb",
  1877 => x"4b7087eb",
  1878 => x"03abb7c0",
  1879 => x"c087f3fd",
  1880 => x"4d2687c2",
  1881 => x"4b264c26",
  1882 => x"00004f26",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00040000",
  1887 => x"ff010000",
  1888 => x"c8f30882",
  1889 => x"50f364f3",
  1890 => x"018101f2",
  1891 => x"ff1e00f4",
  1892 => x"e1c848d0",
  1893 => x"ff487178",
  1894 => x"c47808d4",
  1895 => x"d4ff4866",
  1896 => x"4f267808",
  1897 => x"c44a711e",
  1898 => x"721e4966",
  1899 => x"87deff49",
  1900 => x"c048d0ff",
  1901 => x"262678e0",
  1902 => x"1e731e4f",
  1903 => x"66c84b71",
  1904 => x"4a731e49",
  1905 => x"49a2e0c1",
  1906 => x"2687d9ff",
  1907 => x"4d2687c4",
  1908 => x"4b264c26",
  1909 => x"ff1e4f26",
  1910 => x"ffc34ad4",
  1911 => x"48d0ff7a",
  1912 => x"de78e1c0",
  1913 => x"faebc27a",
  1914 => x"48497abf",
  1915 => x"7a7028c8",
  1916 => x"28d04871",
  1917 => x"48717a70",
  1918 => x"7a7028d8",
  1919 => x"c048d0ff",
  1920 => x"4f2678e0",
  1921 => x"48d0ff1e",
  1922 => x"7178c9c8",
  1923 => x"08d4ff48",
  1924 => x"1e4f2678",
  1925 => x"eb494a71",
  1926 => x"48d0ff87",
  1927 => x"4f2678c8",
  1928 => x"711e731e",
  1929 => x"caecc24b",
  1930 => x"87c302bf",
  1931 => x"ff87ebc2",
  1932 => x"c9c848d0",
  1933 => x"c0487378",
  1934 => x"d4ffb0e0",
  1935 => x"ebc27808",
  1936 => x"78c048fe",
  1937 => x"c50266c8",
  1938 => x"49ffc387",
  1939 => x"49c087c2",
  1940 => x"59c6ecc2",
  1941 => x"c60266cc",
  1942 => x"d5d5c587",
  1943 => x"cf87c44a",
  1944 => x"c24affff",
  1945 => x"c25acaec",
  1946 => x"c148caec",
  1947 => x"2687c478",
  1948 => x"264c264d",
  1949 => x"0e4f264b",
  1950 => x"5d5c5b5e",
  1951 => x"c24a710e",
  1952 => x"4cbfc6ec",
  1953 => x"cb029a72",
  1954 => x"91c84987",
  1955 => x"4bd6f8c1",
  1956 => x"87c48371",
  1957 => x"4bd6fcc1",
  1958 => x"49134dc0",
  1959 => x"ecc29974",
  1960 => x"7148bfc2",
  1961 => x"08d4ffb8",
  1962 => x"2cb7c178",
  1963 => x"adb7c885",
  1964 => x"c287e704",
  1965 => x"48bffeeb",
  1966 => x"ecc280c8",
  1967 => x"eefe58c2",
  1968 => x"1e731e87",
  1969 => x"4a134b71",
  1970 => x"87cb029a",
  1971 => x"e6fe4972",
  1972 => x"9a4a1387",
  1973 => x"fe87f505",
  1974 => x"c21e87d9",
  1975 => x"49bffeeb",
  1976 => x"48feebc2",
  1977 => x"c478a1c1",
  1978 => x"03a9b7c0",
  1979 => x"d4ff87db",
  1980 => x"c2ecc248",
  1981 => x"ebc278bf",
  1982 => x"c249bffe",
  1983 => x"c148feeb",
  1984 => x"c0c478a1",
  1985 => x"e504a9b7",
  1986 => x"48d0ff87",
  1987 => x"ecc278c8",
  1988 => x"78c048ca",
  1989 => x"00004f26",
  1990 => x"00000000",
  1991 => x"00000000",
  1992 => x"005f5f00",
  1993 => x"03000000",
  1994 => x"03030003",
  1995 => x"7f140000",
  1996 => x"7f7f147f",
  1997 => x"24000014",
  1998 => x"3a6b6b2e",
  1999 => x"6a4c0012",
  2000 => x"566c1836",
  2001 => x"7e300032",
  2002 => x"3a77594f",
  2003 => x"00004068",
  2004 => x"00030704",
  2005 => x"00000000",
  2006 => x"41633e1c",
  2007 => x"00000000",
  2008 => x"1c3e6341",
  2009 => x"2a080000",
  2010 => x"3e1c1c3e",
  2011 => x"0800082a",
  2012 => x"083e3e08",
  2013 => x"00000008",
  2014 => x"0060e080",
  2015 => x"08000000",
  2016 => x"08080808",
  2017 => x"00000008",
  2018 => x"00606000",
  2019 => x"60400000",
  2020 => x"060c1830",
  2021 => x"3e000103",
  2022 => x"7f4d597f",
  2023 => x"0400003e",
  2024 => x"007f7f06",
  2025 => x"42000000",
  2026 => x"4f597163",
  2027 => x"22000046",
  2028 => x"7f494963",
  2029 => x"1c180036",
  2030 => x"7f7f1316",
  2031 => x"27000010",
  2032 => x"7d454567",
  2033 => x"3c000039",
  2034 => x"79494b7e",
  2035 => x"01000030",
  2036 => x"0f797101",
  2037 => x"36000007",
  2038 => x"7f49497f",
  2039 => x"06000036",
  2040 => x"3f69494f",
  2041 => x"0000001e",
  2042 => x"00666600",
  2043 => x"00000000",
  2044 => x"0066e680",
  2045 => x"08000000",
  2046 => x"22141408",
  2047 => x"14000022",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
