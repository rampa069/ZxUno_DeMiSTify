library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"14141414",
     1 => x"22000014",
     2 => x"08141422",
     3 => x"02000008",
     4 => x"0f595103",
     5 => x"7f3e0006",
     6 => x"1f555d41",
     7 => x"7e00001e",
     8 => x"7f09097f",
     9 => x"7f00007e",
    10 => x"7f49497f",
    11 => x"1c000036",
    12 => x"4141633e",
    13 => x"7f000041",
    14 => x"3e63417f",
    15 => x"7f00001c",
    16 => x"4149497f",
    17 => x"7f000041",
    18 => x"0109097f",
    19 => x"3e000001",
    20 => x"7b49417f",
    21 => x"7f00007a",
    22 => x"7f08087f",
    23 => x"0000007f",
    24 => x"417f7f41",
    25 => x"20000000",
    26 => x"7f404060",
    27 => x"7f7f003f",
    28 => x"63361c08",
    29 => x"7f000041",
    30 => x"4040407f",
    31 => x"7f7f0040",
    32 => x"7f060c06",
    33 => x"7f7f007f",
    34 => x"7f180c06",
    35 => x"3e00007f",
    36 => x"7f41417f",
    37 => x"7f00003e",
    38 => x"0f09097f",
    39 => x"7f3e0006",
    40 => x"7e7f6141",
    41 => x"7f000040",
    42 => x"7f19097f",
    43 => x"26000066",
    44 => x"7b594d6f",
    45 => x"01000032",
    46 => x"017f7f01",
    47 => x"3f000001",
    48 => x"7f40407f",
    49 => x"0f00003f",
    50 => x"3f70703f",
    51 => x"7f7f000f",
    52 => x"7f301830",
    53 => x"6341007f",
    54 => x"361c1c36",
    55 => x"03014163",
    56 => x"067c7c06",
    57 => x"71610103",
    58 => x"43474d59",
    59 => x"00000041",
    60 => x"41417f7f",
    61 => x"03010000",
    62 => x"30180c06",
    63 => x"00004060",
    64 => x"7f7f4141",
    65 => x"0c080000",
    66 => x"0c060306",
    67 => x"80800008",
    68 => x"80808080",
    69 => x"00000080",
    70 => x"04070300",
    71 => x"20000000",
    72 => x"7c545474",
    73 => x"7f000078",
    74 => x"7c44447f",
    75 => x"38000038",
    76 => x"4444447c",
    77 => x"38000000",
    78 => x"7f44447c",
    79 => x"3800007f",
    80 => x"5c54547c",
    81 => x"04000018",
    82 => x"05057f7e",
    83 => x"18000000",
    84 => x"fca4a4bc",
    85 => x"7f00007c",
    86 => x"7c04047f",
    87 => x"00000078",
    88 => x"407d3d00",
    89 => x"80000000",
    90 => x"7dfd8080",
    91 => x"7f000000",
    92 => x"6c38107f",
    93 => x"00000044",
    94 => x"407f3f00",
    95 => x"7c7c0000",
    96 => x"7c0c180c",
    97 => x"7c000078",
    98 => x"7c04047c",
    99 => x"38000078",
   100 => x"7c44447c",
   101 => x"fc000038",
   102 => x"3c2424fc",
   103 => x"18000018",
   104 => x"fc24243c",
   105 => x"7c0000fc",
   106 => x"0c04047c",
   107 => x"48000008",
   108 => x"7454545c",
   109 => x"04000020",
   110 => x"44447f3f",
   111 => x"3c000000",
   112 => x"7c40407c",
   113 => x"1c00007c",
   114 => x"3c60603c",
   115 => x"7c3c001c",
   116 => x"7c603060",
   117 => x"6c44003c",
   118 => x"6c381038",
   119 => x"1c000044",
   120 => x"3c60e0bc",
   121 => x"4400001c",
   122 => x"4c5c7464",
   123 => x"08000044",
   124 => x"41773e08",
   125 => x"00000041",
   126 => x"007f7f00",
   127 => x"41000000",
   128 => x"083e7741",
   129 => x"01020008",
   130 => x"02020301",
   131 => x"7f7f0001",
   132 => x"7f7f7f7f",
   133 => x"0808007f",
   134 => x"3e3e1c1c",
   135 => x"7f7f7f7f",
   136 => x"1c1c3e3e",
   137 => x"10000808",
   138 => x"187c7c18",
   139 => x"10000010",
   140 => x"307c7c30",
   141 => x"30100010",
   142 => x"1e786060",
   143 => x"66420006",
   144 => x"663c183c",
   145 => x"38780042",
   146 => x"6cc6c26a",
   147 => x"00600038",
   148 => x"00006000",
   149 => x"5e0e0060",
   150 => x"0e5d5c5b",
   151 => x"c24c711e",
   152 => x"4dbfdbec",
   153 => x"1ec04bc0",
   154 => x"c702ab74",
   155 => x"48a6c487",
   156 => x"87c578c0",
   157 => x"c148a6c4",
   158 => x"1e66c478",
   159 => x"dfee4973",
   160 => x"c086c887",
   161 => x"eeef49e0",
   162 => x"4aa5c487",
   163 => x"f0f0496a",
   164 => x"87c6f187",
   165 => x"83c185cb",
   166 => x"04abb7c8",
   167 => x"2687c7ff",
   168 => x"4c264d26",
   169 => x"4f264b26",
   170 => x"c24a711e",
   171 => x"c25adfec",
   172 => x"c748dfec",
   173 => x"ddfe4978",
   174 => x"1e4f2687",
   175 => x"4a711e73",
   176 => x"03aab7c0",
   177 => x"d9c287d3",
   178 => x"c405bfc7",
   179 => x"c24bc187",
   180 => x"c24bc087",
   181 => x"c45bcbd9",
   182 => x"cbd9c287",
   183 => x"c7d9c25a",
   184 => x"9ac14abf",
   185 => x"49a2c0c1",
   186 => x"fc87e8ec",
   187 => x"c7d9c248",
   188 => x"effe78bf",
   189 => x"4a711e87",
   190 => x"721e66c4",
   191 => x"87f9ea49",
   192 => x"1e4f2626",
   193 => x"c348d4ff",
   194 => x"d0ff78ff",
   195 => x"78e1c048",
   196 => x"c148d4ff",
   197 => x"c4487178",
   198 => x"08d4ff30",
   199 => x"48d0ff78",
   200 => x"2678e0c0",
   201 => x"d9c21e4f",
   202 => x"ff49bfc7",
   203 => x"c287eadf",
   204 => x"e848d3ec",
   205 => x"ecc278bf",
   206 => x"bfec48cf",
   207 => x"d3ecc278",
   208 => x"c3494abf",
   209 => x"b7c899ff",
   210 => x"7148722a",
   211 => x"dbecc2b0",
   212 => x"0e4f2658",
   213 => x"5d5c5b5e",
   214 => x"ff4b710e",
   215 => x"ecc287c7",
   216 => x"50c048ce",
   217 => x"dfff4973",
   218 => x"497087cf",
   219 => x"cb9cc24c",
   220 => x"dacb49ee",
   221 => x"c24d7087",
   222 => x"bf97ceec",
   223 => x"87e4c105",
   224 => x"c24966d0",
   225 => x"99bfd7ec",
   226 => x"d487d705",
   227 => x"ecc24966",
   228 => x"0599bfcf",
   229 => x"497387cc",
   230 => x"87dddeff",
   231 => x"c1029870",
   232 => x"4cc187c2",
   233 => x"7587fefd",
   234 => x"87efca49",
   235 => x"c6029870",
   236 => x"ceecc287",
   237 => x"c250c148",
   238 => x"bf97ceec",
   239 => x"87e4c005",
   240 => x"bfd7ecc2",
   241 => x"9966d049",
   242 => x"87d6ff05",
   243 => x"bfcfecc2",
   244 => x"9966d449",
   245 => x"87caff05",
   246 => x"ddff4973",
   247 => x"987087db",
   248 => x"87fefe05",
   249 => x"f7fa4874",
   250 => x"5b5e0e87",
   251 => x"f80e5d5c",
   252 => x"4c4dc086",
   253 => x"c47ebfec",
   254 => x"ecc248a6",
   255 => x"c178bfdb",
   256 => x"c71ec01e",
   257 => x"87cbfd49",
   258 => x"987086c8",
   259 => x"ff87ce02",
   260 => x"87e7fa49",
   261 => x"ff49dac1",
   262 => x"c187dedc",
   263 => x"ceecc24d",
   264 => x"cf02bf97",
   265 => x"ffd8c287",
   266 => x"b9c149bf",
   267 => x"59c3d9c2",
   268 => x"87cffb71",
   269 => x"bfd3ecc2",
   270 => x"c7d9c24b",
   271 => x"ebc005bf",
   272 => x"49fdc387",
   273 => x"87f1dbff",
   274 => x"ff49fac3",
   275 => x"7387eadb",
   276 => x"99ffc349",
   277 => x"49c01e71",
   278 => x"7387dafa",
   279 => x"29b7c849",
   280 => x"49c11e71",
   281 => x"c887cefa",
   282 => x"87fdc586",
   283 => x"bfd7ecc2",
   284 => x"dd029b4b",
   285 => x"c3d9c287",
   286 => x"dec749bf",
   287 => x"05987087",
   288 => x"4bc087c4",
   289 => x"e0c287d2",
   290 => x"87c3c749",
   291 => x"58c7d9c2",
   292 => x"d9c287c6",
   293 => x"78c048c3",
   294 => x"99c24973",
   295 => x"c387cf05",
   296 => x"daff49eb",
   297 => x"497087d3",
   298 => x"c00299c2",
   299 => x"4cfb87c2",
   300 => x"99c14973",
   301 => x"c387cf05",
   302 => x"d9ff49f4",
   303 => x"497087fb",
   304 => x"c00299c2",
   305 => x"4cfa87c2",
   306 => x"99c84973",
   307 => x"c387ce05",
   308 => x"d9ff49f5",
   309 => x"497087e3",
   310 => x"d60299c2",
   311 => x"dfecc287",
   312 => x"cac002bf",
   313 => x"88c14887",
   314 => x"58e3ecc2",
   315 => x"ff87c2c0",
   316 => x"734dc14c",
   317 => x"0599c449",
   318 => x"c387cec0",
   319 => x"d8ff49f2",
   320 => x"497087f7",
   321 => x"dc0299c2",
   322 => x"dfecc287",
   323 => x"c7487ebf",
   324 => x"c003a8b7",
   325 => x"486e87cb",
   326 => x"ecc280c1",
   327 => x"c2c058e3",
   328 => x"c14cfe87",
   329 => x"49fdc34d",
   330 => x"87cdd8ff",
   331 => x"99c24970",
   332 => x"87d5c002",
   333 => x"bfdfecc2",
   334 => x"87c9c002",
   335 => x"48dfecc2",
   336 => x"c2c078c0",
   337 => x"c14cfd87",
   338 => x"49fac34d",
   339 => x"87e9d7ff",
   340 => x"99c24970",
   341 => x"87d9c002",
   342 => x"bfdfecc2",
   343 => x"a8b7c748",
   344 => x"87c9c003",
   345 => x"48dfecc2",
   346 => x"c2c078c7",
   347 => x"c14cfc87",
   348 => x"acb7c04d",
   349 => x"87d3c003",
   350 => x"c14866c4",
   351 => x"7e7080d8",
   352 => x"c002bf6e",
   353 => x"744b87c5",
   354 => x"c00f7349",
   355 => x"1ef0c31e",
   356 => x"f649dac1",
   357 => x"86c887fd",
   358 => x"c0029870",
   359 => x"ecc287d8",
   360 => x"6e7ebfdf",
   361 => x"c491cb49",
   362 => x"82714a66",
   363 => x"c5c0026a",
   364 => x"496e4b87",
   365 => x"9d750f73",
   366 => x"87c8c002",
   367 => x"bfdfecc2",
   368 => x"87d2f249",
   369 => x"bfcbd9c2",
   370 => x"87ddc002",
   371 => x"87cbc249",
   372 => x"c0029870",
   373 => x"ecc287d3",
   374 => x"f149bfdf",
   375 => x"49c087f8",
   376 => x"c287d8f3",
   377 => x"c048cbd9",
   378 => x"f28ef878",
   379 => x"5e0e87f2",
   380 => x"0e5d5c5b",
   381 => x"c24c711e",
   382 => x"49bfdbec",
   383 => x"4da1cdc1",
   384 => x"6981d1c1",
   385 => x"029c747e",
   386 => x"a5c487cf",
   387 => x"c27b744b",
   388 => x"49bfdbec",
   389 => x"6e87d1f2",
   390 => x"059c747b",
   391 => x"4bc087c4",
   392 => x"4bc187c2",
   393 => x"d2f24973",
   394 => x"0266d487",
   395 => x"de4987c7",
   396 => x"c24a7087",
   397 => x"c24ac087",
   398 => x"265acfd9",
   399 => x"0087e1f1",
   400 => x"00000000",
   401 => x"00000000",
   402 => x"00000000",
   403 => x"1e000000",
   404 => x"c8ff4a71",
   405 => x"a17249bf",
   406 => x"1e4f2648",
   407 => x"89bfc8ff",
   408 => x"c0c0c0fe",
   409 => x"01a9c0c0",
   410 => x"4ac087c4",
   411 => x"4ac187c2",
   412 => x"4f264872",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
